PK   상V|�">8  -@    cirkitFile.json�}�n%7��4��.��a�Lֿv����1�Y�6��F�j$U���h_f�i�<R�N^�a���T�v͠-)����`|���������ۻ~����������ˋ�����_���۫�����/w���.���~/~|��]_w�m,�SD��;S4me
�uS4u��v>P��z�v�����^�/��Ԏ���N�1p%��ac�JP;�����v���+A�J6���Q����ooo���]W;���Cma��E��(HYo;E�%�<���b��+AE-<W�����⮾��Evoo�뻫����/L���T��Ĭ |=�j��5����6E��Q����ֈ?��a��(�C[DD�|�""
���Qp� ⋈(��[DD�u���T~����8�F��!��Fq4dր�wG�׀��}6[DD��p�)����|�w�l�g7�#��>tŭQ�� �?i�P��v�?�ED���-"��El`������Q��x㘎�8�+�5�l�ִVi�5��	�������"b�ÚN��C���w�l���^uhl��
�P(��Z��<�j�U���K�����$���%��w���@,��ysn�c�I{�9-�d�g�Pˍ�Հ�9@Ѿ�L��Gi����?ҲED���-B��-�ED�ŗ�ѫ��e��ά>o�&�gמ[}���X3iN������5�g\��q�6U8V�-�\6�l���4[DD���""
�8�Q��i�����=Ԯ��l�"�ED�ҙ������F,t�YH��1�8�dtB��NT�2�	Lܾb<=A�]�X�i����N�Vw�;(:¢�<�;��a����;��a������;(:¢S;�՝������Ԯ����������]�����fGx;�7����<Hl�G`|��Xhn�&'`v2={�������fRrl��I�����������4���������T����ҹ$���t����҉*���������Y0���������)6����������;��6��`�_:9���`�_:��zy����?4�`�_:�	��`�_���`�_:$��`�����Eʃ�o��3�5�t˃Q?��L�&���/s|�欘��~4��`�_:�ޟf?X|Ɨ���f?X|Ɨ�ك�f?X|Ɨ����`��af?�~��`���%D@ʃ�o���pe���Q?�<0y��#0����?0y��#0��y�?0���#0��3�?0}��#0����?�/X|Ɨ�����/X|����gs�b�䅭z0���L�X�5l�RJ����	����RF��Чs��s��ɂ��',>Z�w���Ե`�d��	����R*"����	����R%����	����R�'����	����R�*���4a�_J���4a�_�����`�_J����`�_����`�����Bʃ����k>��<g`���-�;�97��S�>X|Ɨ�ҁ��>X|Ƨ��A��>X|��}LW�MuP��S	fNX|Ɨ��fNX|ƗR.��fNX|t���Ӽ�[��O3]n,>͕�9�#/��į��n"�Q+n��wC�j�fvc��9�7�&�|s�Wq��_���Onb>��I���y��<�Cͮ�Z~�}k��%[�3���Zܭ����_4�칖c>��yfvn���W��&�Ξu�:��̾7��u�n̍�,ǭK��O���yָ��C�c���w���.�Z~=�o78ݔ��+��mQ�v(B[S��-5GXEVq�������n#s$/����d@���3o�c~}�f^O'4�g��b������__������Y�ףǬ�ӛZ�_&4���%4�ޣ%4��c%4��#���c}�}U�〬
�u�.��Da&�EE�K�F�^w�H0�U|=(��֍���l�L\?uB��+c`s��Y�׿N�۠����C,���qT�ڦ�m�?����G!�z��hYTF�66cm�+T=t���X�c��*���z�M��1�h��Ǻ���
j�3�B�Q8>��:���L��1��U4wUua�65�d�COmP�ű��Yŏ4�wnrYU���5��^}kz����tǺLV���Gs�u���&��6��!������WG��U|��M5��*��Tu4�ઢ��Pt�T�����泊�ݑ/��VQ���.��eQE
Ml���泊�}0U��/L�!q�PTC��5-�.Խm�Y]N�#V�ڡ�]Y�~p�u]䜵
�T��u�Y]N���+j��i�":�2vؾ�Ί�������)u��Y�ǯ�<��=�����ۻ�7?q�������sQ3��]�$H%/�A���� 	R��b���H1�@�Tb�D Ai�.
�Nn�4�G!�P:	Jw����0�D`r����l6�y����4��u�0�M����s�P��s�(Ij�E a�yo��o�$5.S�0�<8�</�$�q9�	��	�}	&I�������5,�FIR�
?�(���r��`~|/�i���'�GIR���$���LL0?�a~%iL��U4̏�
�j��0?����} :����Q�R�X&�L
n*��GIJ�Aa��ӥ��0L0?n`��^�0���31��q���-�	������0�4NO��`~%iܰ�U,̏[��-J���	7'>z߲2�i��`~���8JҸ��,̏[�GIJɦ`�`~���8JRJ�[���q7z�@�j������{���k̏����u�˖�	��ݣ��{όnus�������ɢGI�x���q�����	��̏�$�l0L�Ӕ��`��%,GIJ�`�V$�O�/z�I�E;c���`��p�`U�i�LkMse ��V��v��p�@�J`%�j7�G�
ԫV�y��^��
1��J"Xc$��iB�$������u���	�$�U�I�R�z��J"X�n��.�W	�$�U�I
�R�z��J�X�`Nb��%�ׁZ�A��6��V�u	�.�E2ċd��Z�T�ڴ�\F�2�K-ɠM{�et+��DВڴ�_F�2,L-ɠMgdt+��DВ�tCF�2lL-ɠMgJdt+��DВ�t6FF�2�L-ɠMg|ddx�Z�A��*��V����%��̕�n�VĄ��dx���eZ����%����nex�Z�A�����V����%��L��nex�Z�A��V��V��-�E�1��MgDet+��D��2Z�����eZ����%��̮��$^&��dЦ��2���e"hIm:C-�[^&��dЦ��2�ڭ(�]Q��^fdx�Z�A�����V��-�Eķ"hS����2�$�6�J�ѭ/AK2hS����2�$�6宐ѭ/AK2hS�Z^&��dЪ�;�����e"h�_��j�/�2�l-"A�r���V����%�)G��n�N�	%��eV��MomC)Af�l-����2+��DВڔ�HF�2�L-ɠM9�dt+��DВڔ�JF�2�L-ɠM9�Dt�dx�Z�A�r���V����%�)Ǚ�nex�Z�A�r���V����%�)県nex�Z�A�r���V(ˇ�z�Zup�/R�2�L��Zc�u2����2�$�6�d�ѭ/AK2hSnI���2�����J^V��2�$�6���ѭ/AK2hS�R���2������]��:[!��%�u�M�);ݻI�%�v�F)+�i7JY�&�Q�J�R�r�Q�[����d��(e%�F)�ҳ;O6Js>�/�ju��ί��*f����z[�`�w�֭bVR�o�rk�V1^�st���4�[ŌV<��e��{t���L����1��y��ъ�3o��ⵋ%���x~7�V1��/��*�ъ��hl3Z��ꋭb��Oo��:�b���?�i-�)
eWX_ۢ��P���.(�[jNG5YR0XNYRN�'��P��}��"��m����]�OzY�G��Щ�(K�����\��S>8K���e��ڍRN�YRN��YRN�YRV�
�ju���C��o�}���1��o��р���ls��X��:]4���ۄ���t������i�%��-��֍���cml�L\?uB�ͮ���i,YRNb!�m�UTj�!Ji}�8�
_m��6۟ƒ%����Zo����FV7Em�+T=t���X��6ʒ��rr�����_�C�^�*���
j�3�B�Q8]�,)'k�%S��c��U�B���vm(jr�3=�AQg�i�dI9��޹!�z�U��X���uѷ�w]��M����������G�69�е���0��t���:�%K�I,M5��*��Tu��UE]��謩t�;�}FeI9�ő/��VQ���.��eQE�M��:������2����&�H@(��j՚�|�޶��#��v�zW�\a]�I�"��m0^�}�e�n���X5M�]�f=C�F�IqP�H�*�X��<���(f�p�����7?}�������pW_?Ƿ��1��}?� 	R�A����$H���$H��$H�|�$H���$H�<�$H���$H��5�E�6�m��6�7J��O#`0�|7��7J��Op`0��7�8J��/�a0�|8��8J��/b0�����q�$�_��`��߸ ��5̏�$��,̏k�GIR��a&��0?������L0?�a~%I�W�1t��̏�$�\�0L���T
̏�GIJ9a�`~���8JR�Q�����Q�RN4&��0?���rp�0�����q����	�	7'����q��(I)7̏[�GIJ�``�`~���8JR�=[���q��(I)�̏;�GIJ�`�p����M�w0?������0�����q��t��	��K�GIJg|a�`~����5I����΃������V��v���h�@�J`%�j7;��
ԫV��v��\h�@�J`%��w��u���	�$�5�A"z���h@+�`�1��^g� ��J"X�n��-�W	�$�U�fy��R�z��J"X�n��-�W	�$�5�	�!2�K-ɠM{�et+ĺ�h��"�E2�K-ɠM{�et+þDВڴg^F�2L-ɠM{�et+��DВ�t�AF�2LL-ɠMg1dt+��DВ�t�DF�2�L-ɠMgcdt+��DВ�t�GfaA����%�鬒�nex�Z�A��\��VhELhIL��i^�ex�Z�A�����V����%��,��nex�Z�A��$��V����%��l��nex�Z�A�Έ��V����%�鬫�nex�Z�A����lL��e"hIm:{,�[^&��dЦ3�2���e"hIm:.�[�݊B�ex���eF����%��l��nex�Z�A�r��V����%�)W��nex�Z�A�r>��V����%�)w��nex�Z�A�rp�����2�$�6��ѭ/AK2hSN���2�$�6�v�ѭ/AK2hS��
�$:J&�ˬ/�2�L-ɠM9�dt+��DВڔ�HF�2�L-ɠM9�dt+��DВڔ�JF�2�L-ɠM9�Dt�dx�Z�A�r���V����%�)Ǚ�nex�Z�A�r���V����%�)県nex�Z�A�r���V(ˇP�^�dx���e"hIm�e(�[^&��dЦ��2���e"hIm�-)�[^&��dЦ�"�-ex�Z�A�r}��V����%�)g��nex�Z�C���vVw�-��鋺�&]��m�ȷd��a�(e%7�F)+�d7JY��Q�J��RVreo����z���|���d��(e%��V�/�z�.}�*c�kW�n���L������5�[�`�Xc�x��̭b0V�vK�V1+^�r���ݸ�UƊ��5�:�b�x���b��N7eA��
�k[T������tK��&K
���%�d�^uhl��
�P(�����<�j�UyZ/YRN�%K�I�dI��夛ɒr��dI9�d����1YRN��,)'=L�Ձ�c����<1�=��9i�V�N�`��6�/**]b��|�;s��dI9�NeYٺ1�0}����)�뇢�B��ٕqx9�%K�I,����J�?D)�/GU᫡m�ކ`��X����\����2��ꦨMp���Ζ]���FYR0XNw%�jg�/ڡ�Q/FM�w5�K��(d�m9RN{�)���Ch�W��r�۵��ɥ�4��E�u���%�tK{��QVU��c���Eߚ�u�G7]Fo̒rK�B��b����B�Fg7��4C�Qӓ��4�,)'�4�ڪ�SձWu����ҍ���m�%�$G��*[D}�Қ�ڗE�/4�
�6ʒr�`�6z\_��C"����-TkZ�]�{�f�n��Ӷ�ڡ�]Y�~p�u]�&�
�T��u_w��#�$EM�CWD�YF�з�cR��*���rJe`ɒ��ϗ�ǿ�J�^����]����⇫��~�����iwu�������7_�᛬p��KƷ+^�������o�����m�bT�O;���d��Ő��;@®JG3d/�Z3$g�7��qj!��\u���",%L��p�0�czb���NϺ�g/���Cn$9�z�W�+��G�}�kxG��G	QDn ī�j���>�s�d�����[����N��������|>�?o_�󬶯X��qR�^�c~���.��\��Y��W:]f�,i�Ú�u��1����PJQ-�-S`��Fά09�1$gy\���,��岰L%�TC���Mȿf�W�4L��+K�\8P�	嘹�����¶ݖ��u���r�L�n?eM�0C��,�v	��"0�4;�<\q;��TP�.��"ͥ8l[�N��<�͚LׅRF���*vsp�Μf��9n?���<g��yV��S�1�=ö�3ᜏ��xB�YK<�	��	�SqPUm?R��<sV<��g2Jl��{�}�mu��׾��7��Ϋ�#�����_p� w w3 wO skx���oT[ �i�W~:����>]u!\0x�����7mŗ�h8�Vģ^dG"zc"`�W܎��]rn�㯠�Fc����k�������Z���&Vns����.^`G-�U��\u�2
��^�"��ر���c�L��Fěd��혐v!�v�
��;���bc< `< `�< `�<�:����a��rw�cPp7�Z��"�S�@��p� ��G�  '�:�<�0#��Qz�X!�N# �3�� S^\�9�e_�@-�(=c��EΎ`z�	�|��e-�~�J �x�[?>�S(��l�a����"gR���GS ;�O�X:'!q�T��?Im�2���a.^�4{w(;�A����|DJnq:{�=���2�<"xy�"�nG� @�'�0������	�)���;O��w��~̑�l�>R[��Om����'M1�y��7��N�}��'؇`?�Y؊�"�� ނ�?P��y:����	�I�3�O�@�4*��橅A�6�+�pc[ȠB�-�\8�$����~���=�~���ˋ��wW7�������x����a؋�=���]uo~�M���x��������-B�?1Q�E���(&
�5^��D���K�(�"�x�#[�/�T����|P_5lj���P5ܓZ��Լ�X'
i/�����LX �;^�9����e���\ �L �̗��w�sq �2�}(dD G̗�ҾB>��Հ��/C�u{>Dh��m�.Z3w�k�{eL`1W�4���e���Ӫ)�5ڋ��8_��q}z3�V�i/����bΨh�k� �̗�-�5�eD �̗q \3_Fā�x ���|�2T�K��;p�<al Η/C�I^>����=GX�@�/#� x[��q��LŬM?�Ʌp�|��Y�ŜU� _l�1�b�YĤ��G6ܔH Om��/c�N��-�S[���ˈ8 ��/#� �f��s�@�/cL�33[���H.���t6��݂kf�����5+���Era-�`0���Hv�@L͗q <5_F���|*����XXd�(��/#� �|`c.�}|�%X�g��g~��)_�,�;���=�-i
�%����� �7D�?,>�S;֟�����")�ς���G`|1T�ρ���G`|1� �������΃������#0>���������#0>�<�D�?,�Y"���O�gl�O��n �EHh�i�+Z�pRg%hZ2M�����73�X��-�h���
!����h��
!����h�9!���D�y�<w��h�Bh�FHh�i�?Z�h�FHh���Z�hFHh���zM[�	�P�2�Bbt��-`�j�S*�C��
��h4O�h�FHh�� Z�h�FHh��Z�h�FHh���Z�h�FHh�j��*����Ts�
�:H[�Q)����3�?)x��,F�Y!�����$hFHh��t%Z�hFHh��d(Z�hFHh��T+Z��a�ahc�,ƠY!��Y�G�@�g'[�������h��I!��S�h�I!��#�h�Y!����h�i!����`Z4m#$4BupU+F�h�F8��vv2���J��/��b�'`����C�U�&5`��F�rY�u?�?�&5Mj���^��#��߲nL9D�*E�0BB#L	O�:D�0BB#L�Z�:D�0BB#L�f�:D�0BB#LIr�:thRFHh�)�Z�hRFHh�)Z�hFHh�)uZ�h�FHh�)�Z�h�FHh�))Z����'�b���2h�U��-`���p�F��4�qhFHh�)�Z�hFHh����<��,�p~/��r�5P�IM�&5`��F��ߡu�&5`��F���u�&5`�t
���:gI�^��,?K����,������9��/$�-�fY7��eR�X~~��]�}���W���i�����a�*�k��{��
�%@�*`�T~� �	���*`��w���U�77��$�[�������8�_s�<��/"�~��[Z��[�&��(�S,��mź�{����/��*�H��6np�)
eWX_ۢ��P���.D�-5��������R���-��Ua
E0Q�>t�'[�*w.h��g�[�ae`��poC�g��w����q�se�;uC�FqG�۬�G�۬�GF۬��[Mq��W|s����X��5�k�9O�ܺ�|s���k8V��<y�]���U����E3���M苊J���!�;s�sg�?�˲�ucla�X[;S�E݅)�+�@t��Y�|���AWQ��X��E�*|5�M��l��Y反\��V}�P�[��	�P��ٲ�ce��?�<��GFNoZ��E;4>�ߨ�i����:c)T�c�����U�����?�FyM_�C]خEM.u���6(�;V������;7�����X��J�U���5��b�k���'����Gӷu��&�6��!������WǾ�U����jmUօ��h��UE]��謩t�;��Q�g�?�}G��*[D},ߚ�ڗE-)4�m����*�������|a�)`E5Tm�ZӒ�B������?f��ޕE�WX�E�P���N��x]�uw��r������}�+�+c����(]��rJ�~V������P��=�����7?]���7__� &)XHr
:�@��+H|���Xy�pǙ�q�W��DcF�1C�8�7N<�Tb�(���9����H�ǥ�qBA�:�0�D$u��jeП9�X0'A�;~.'���X ':8(�3��?5�Ԗ1�,�;g�8����
���9��@��;(��+��S
�8�g�#x���7�C����0�9�7Z�����ɺ)kyn"k^Q{Pѳn@�Py֬�%�v�0Lm8֬!G���Ϋ���ac�.�Bu�[ּg7����hnu8�^ks
�����8nuX�&vQ��m,�����څ�!*sƘ�<��"���{f�;/�3G��ͺ�#����t��j����Ӝ艩��66T����p����o�y����%�7��z���ޑ:�Kf�0p��i�Hs�l�,��:n ����	7�K.B�CӴ��6憺�cu����)Y9g�^ 7���R�o���I�x��ih!�ч�2&a'P8ܒt���y�a�|�7d�r��=d�x�~>�����aw]7�u�I;ę��.��?�J��G��?2�����z|�������Gz��=>r�G��j�(<>
�G���=����{�Os���+�+��TLs���h�{O��y��S��B��tIseғ%����Z�\-�}��뮟����x4o=��=׋~����A?�A/��I���7���ݳ^yu3���I�.Z������]��o�����U�����u?<���/������w�C�����/�n��wW�����ۛ���n����nҬ�M�}�==���k}�.�����2����U������/n~�^����>>���������������wWw}w��!�#6���ͻ�n���w� <�������- I�Gϫ��ۨ��_U��}���2��Em&����.��g�)�s��V�E�b�U�����qj������i�e��1//n�bs�{0���?�Ww�u�؀_��ݥ�"�6�g�x��9���A�Wصf���P+%J��z����v��^+A+%\X)Q����_��'���z��W夾O<�<pk%�Z	�Vb���e5��ӃY+<=���ӃY+<=���ӃY+<>��Bz0��.�eg�������.�f���\�����?����o..����ƿ8R�,�2��/�^�	�+}Sն�����^�F��/�_���lת�j*U�¶�/j3P���k�n�Ʋ����Y���WU�ir�>�󴠬�N�u���ߗ����w�
�un膢7i����t�t����T�+x���퓈?F�|��>���]]w�$۔>*z��QrtDu�uј����ֽT������ዷ��3)a Uj]M�5�PT��������߂��^�����(�{�,�����vUAՠMe����X�������S��~���+�,����gs3J�~��OOf���_��?}���/o�~�uw������/�2j�r����u,�ܸbmc�辠�T��L�zlm�����ݫ5����&���mZ�b�V����0����aɸ�(W�J�0�/�C_�ب>��5�Tͪq��e�����*vMYT];G�M�ԅ�=n\���o.�z{ս��޽�����O�|s���?�ӫ��W?޾��?y��~�]�_�z�}u����m��ķ������(���vY����͂���m_?����υ��_���{s��R]^�������Mdl�����2znS^��cu��Y����h�W_=��n��������^�h0����SAΕ����z[�����n�!��!H�7e����S�84*�ʃ8�j{P}Tp��(�ܪ�!P]_�]���~'e헚�I��7�HIW��č��ޏGZ�����y�Ҿ�1�MO^GJ\�����8V�>Ix|��N�o�͌*��7q��{w����7ݻT���ۚI���*E��?;�kg�U�m���\�U_�f(�W�HǱL�A�n����Y�����v�e������
)�2F鑒W��_�gO����&��澆��~��}z��>>p�^��x�>=�D���i��M�)#x��C�PV�����g���x���?����D.�	t���n�.VO{Me��5�/}d4�������T��ϣ�n��a*ň�-c8���kK=Ζt�����>�]�n�:u���|,#��g����?����K���P�ee�K�,��첦�ЍE�P�u��A�5M�j)Y���,e��p�p�+Jr��6���_� a\�{i��⿫��D�^keȆ�	�Q�����gzy��DY�.�žp�Iu燢luS�}GA�����"��m�y�c2E����L�8�r��q��!R��kz�5q#���_��}������?|��'`k��o���o��$�m.�^���\��*��u��!�Gn7��J�01.),�>�����[�fn(�P@F�&1P�,�ܐ��a�V�����J�ey���_���ٻ�w�q�7����7�V�};���;i�q�fҨcɫ�_뛿�S�2r5]�v��x!PZ����u7E?��G<��`��S��MMs?������k��g�m�Y������1��,鬇����M����g�Mw���g(@��؎Y�?�d�e�f��x�Ξ�iк6������]��k}[���v���$y]�-����A�����F�&�c�@�q�6�<S����h���?��S���ڽ��N��o���#�8h�6F�����|lA?�eA�v1��ch��N�����#�Y��9d��,���o9��8��sa�qx?�u871���:��C�Sww�|6x�~N��-����^�
�m�@tdA�[�Z)��k+eC�5�C�#��̜F��O~��+.h4�gN�_z~�uZ?gÖ�hFD�YL��'����s���DMۖ>����zS���Ƙ�h����ԙ>���l�2+aB�҇�-}��҇�-}���~��O�e���JWƛ���c�Yy<r�ۂ�q+��Lљ<�W��EZ��ٿ4C���r�d�|���u��i���m��~�6=!�k ~}$jo.
�A��?�p�=|�^,U�Z�����]z7�E�����6+�����ۺ���>{��˻���������H������]�ލ���!�v�縷.*���˫��݄gg���Dq⌢���BB���Y��۫��/��F�?}��7��×��Wc�t��������N�������޸\z�2j�5{��&�5��Z�������\���dc�N���-��%ژ[{���毭�9k���9ɲ�����Y������]SĿo�@\����n��qM�Q�E���U�O�y3ӛ����m�-`y\���!ܳ_���J��ZE�߯,�F�{�e�_Ƨ��ag۲��i�3��e��1�:�6�8�L}���ԩ�7�#�`B���x4���͸,��閇��[���K6pfnI�'%��W���[v����Y���? ��qhs�@@������2�	/'oU~1xv�e�[١��Kf�VQc�0�5�r��]6��D���r}KYW�l��b��E��A�}����XÜk�dg&;m`�?� ��߲v%��编kԽ���b�����E���ȥ�Y��=s*��83[�h��A 4�?8|�ꕁ_��Z�?hu�>�J�˱ɧͩ��š��=�\ʬ�`�:��*N�羕�[>�||�&GU�Yr8O=�T�yN���#x�3b�[����/U���<ϘV���[�N�Z6�aP:th OA�iѼ�,�9f�9�+��hge:���@!H#,�F��"Ƥ>��7��"^�y3/im_,���XĤ�����[�`������&����V��2kA���!���.�����]�"#��[�f�	�p���r@��G�z+��t�tH�tN�J�[��;_\.����,c�uS��������l/>�Q��s�~N�6g�byCp�k��P>m�^]�i�"�6��g<�������L���9}rkx@"���%�[�[�	Jt��pD:��=l���2�5~�g�����݊���E&>	;�Ik�&>��oit��`?}-�B5�;��&p��l�GR��z	����1�zFO^3�����<�5����zB]F�&�o>�0�o6���)�׀��\�
m��-�r?��%�[M�f�+5�qέ�X�)f������\�;k�T�0�M[1����R,$`8k'�ù��]V���3M��@2_��w,Kӵ�ݲ�.d�͉K8�ksgۧ�y�ї9���J-Ǎ�ͼ��eLSU�9	�".w�(�����MR��J�b0�F+�2&�=3_�5��C�&�����ˍF��Y䳠n��a�����k�^^�/�z-�XDf<v��|�����~�ANe�����;��.��k�2�Yh��(	'z���(!'9|����0�A�k/8�E���Ց�3�5~�:�:ǚ�oe�t�d���df�m�όp־��>ҜՏ����k�:��y����������CwU_�_�I6t?�r����ͻ���������^��۟/~��PK
   상V|�">8  -@                  cirkitFile.jsonPK      =   >8    