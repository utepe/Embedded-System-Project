PK   U�mV�0��)  ��    cirkitFile.json�ko�ȑ�����'���^�����1�^І� Ӄ�na5Ro���lc��f�t+�X�T�1j�i�$����`d�df䗋m���f��n����������{
���m�S��������fw��۶������=����Ϛm_w�m<fc�L[w.k��e��&k������"_o��\������[ ��!1�Ԃ�X1�Ԃ�81�Ԃ�x1�Ԃ�1�Ԃ��b��)�RfS��̦3H-�%O�b��*幒��Rl"R�ӥ�D��'L��H!O�b�B�4�&"�<m�MD
y�����)6�V��)6)�Sl"R :���i�Sl"R�s��D���N��H!ϝb�B�;�&"�<w�MD
y����P�;�&"�<w�MD
y��� �.ϝN�;�&"�<w�MD
y�����)6)�Sl"R�s�؄�xy�����)6)8�=ho�|{���6Ea��j|�W��|CUV��gE��r�e���'�|�S�Ͷ��u2��|����W����wBo�s�woX� ^�z������خ�vq硪�̓볺�����w���<�A��˛/ov�&"E�p���ћ�t��ț;/o��&"�������Nl�l�����$z*r�SAF�Xy;d�,	2sT��˗7�A԰��\~)�|y�D�2I�e+m���m]��^��Mr))6)�m��D����b�B޶�M�M.o[�&"�\J�MD
�k��������HJA��0�Hn��IH������W�Y&>���_��OP:�ҙ����b}�#,��8���wP:��E=�����JGX��_��.`}�#,]��`}�c}�#,��X�X�A�Kg6%�w%�wP:�ҙM��]�����t<��9�u���Y(��x86�hu��`}A`�A`���#0���2�|����`������|<� �?������'L��VX>��T�����G`>���Xy`����k���,��xb�3X`���S����,��x2��/�O`�a��Â����|<�?����������X>��C�����G`>�.	�X`���=���,��x�*�`���#0O�� �,��xZ0�`���#0Oh��?�|���`��GY��Y�����X>���w�����G`>���X`���%���,���X�`���#0�y ��?�|��X�y������Kk���X>:��lm�dK#�V3-�!v=X�������z
�`�����G`>���z�	z�	X�x���`��#|�μ��,�<X4a��ǅk���&,�����`ф�#0�,��|��2GX��h����4��MX>�q�'�����G`>.�X�`���5���K,���H��)��9���6�?X`��߫�I���v	`��#0�4��]�|��bl`������|\F��]�|��x`������|\��?�v���������N�>�����im��� _v{�߈I^�Ė��8�PWŶW5�?���i�ؕ�O+��<|Z�u�C&}H�O�l]˵����Z�k���P^{�0�f+/�=^~�j���^��Z#=}.:���F�lM���������d�/�����[��K�����G7���*{k�_~��&�6yFU�e��}V�vȪ���2ƶԜ�&.<��t��s�8�M֏�����4�/=��+S	Ͼ�&.+��v&��A�A�jœξ�K:|��t�r,�����@J-p��=J-p��9J-p��5J-p��1����o����xS��l�.sU���66B�s':I���e�ͪ΅ؕ�GV��2�+ߵ�kS�ꊤ�|�</}�8��>�_�U������ʐ�nՉ�'�|v2��l�}�!�Y�̊rh���U��gO:���C[x;ĸ�<��D��Bf��yW�+9uߓ�}�X��犬�"^�3�Y軌����:�t�2|��B����x�fw�io�o��H�Q��ſ����W��W�2�bȐỆ!2"�!�cȐ��1�d�p�C2d��!2ܳ��"�!3�P��em\چ�m�%n�%3�,w,y�,�Q耘`��`	eɌ߲@L�N�$��d�on &X��<��dƯs &\����q��(Kf�2	b��q��(Kf��
b��q��(Kf��
b��q��(Kf�*��<�`ye�+poRp�R`y���8�W��1���q�%�nc��q��(K\������Q��Z�	����}�����~̾�`l�	�p���웗�s��	��=,��,�#QFK�uʘ`y���8�1�1���q�%.�����a̾u�� ���!�]�L�<��ץ�[!,����[�E/d�}��ok˶�L�<`�q�%�|c��� ��(K<I���9,��,�d^,���*K���'�����}�dVg�F!��y�V�����ܭ�p�URa%V���	�[�U��TX�fZ�
n�WVRa��Ků�*Xh��
k���uZ�VRa�}�N�fa<��J*�f3���
��+���ʹF�*Я���j6��Yp�@�j��
+�	��T��*��C�c�u|����d���"�E:�K��thy���ouԗ
-���y��(0Zҡ��:��Qa*��C�st|���ThI���b��VG��В-�)��"S�%Z���[U�BK:�<�G�Â�.S�%Z����[]�BK:�<�JǷJ_Ĕ>���2��ˬ�.S�%Z���[]�BK:�<�OǷ:�L��thyN��out�
-����J���2Zҡ�9�:���e*��C�s]u|���ThI�����L��e*��C�s�u|���ThI���P��VG��В-����hE��:����2���ThI������VG��В-���.S�%Z����[]�BK:�\�AǷ:�L��th�v��out�
-��r�z]�BK:��`�out�
�|�Ѭ|^���e^G��ELyT���.:���e*��C�5jt|�4�Li*��.�:�l���	:��(- ���2���ThI��k��VG��В-�p��.S�%Z�E��[]�BK:�\SKŷAG��В-���.S�%Z�q��[]�BK:�\�MǷ:�L��th�朎out�
-��r�<�*U�P*��,��鲥('�貣�r�ttY��e*��C�5u|���ThI��kK��VG��В-��T�m���ThI��k}��VG��В-�,��.S��4��5��:x�u>���<�>�{�_��Pђ_Z�y���ڴ+�,T�]ie���J+��GΕV���J+խWZY�G���B�Vj>��:P�b�wi�׵f0񻴴�Z3��ך���Қ�k�`�x���|���Y�!��˙�5���(^Z�r�L/������E9֚y���:k͌Q<_�b���\<]�bm����K�>�i�0��Uy����Y��!�ښ���Rs�W�d�r��J�r�y*
;�U㳾*L����EoU7������_��#IV�\�(����
\+��s98Ɋ��%�K�IV�6�IVζ�IV�6�IV���ҢΜ˾if�\�M3c�e�43�\�M33�|y��f��o�"t�͚����>+)�TG������d�|�-�:�E�U��A����3�+ߵ�kS&�)Vβ�y������ѳ�.�B?duWUQÇ<6u�Y���e!S�ʖ�����Ț@eV�C����*ߟgI�r����v賆�xE�6Y��z�|�����%�
��lk]��犬�"�ř�i�.���*;��_Q���W�dsE/���f6���ݮ���<�]��ꦿ�m��|�W#2��!D Cf��"�!3��dȌ}8Ȑ��"�!3�-!D Cf�B�@��������!2��8&E�6.m��6�7ʒ�K,w,y�,���0��7�8ʒٿ��0�r8��8ʒ�.�0���q�%����a���qpX��<��d��k0L�<naye��$a�`y���8ʒ���0���q�%������<�`ye�����poRp�R`y���8���1���q�%�gc��q��(K\?	�����Q��^�	��=,��,q}�8�8,�{XGY�:0&X��<���u#`L�<�aye���>���x��q�%�c��� ��(K<Ƅ�����	����Q�x�,�	��,��,��L,��<����aL�<�������s�fsG�V�S� VI��TX�f6om�WVRa5�ٜQ�U�_5XI��lfu|�V�~�`%֨�T�:+��+���~��_g�{ �`%��GQ��t����j6��=h�@�j��
���j������J*�f3�׃�
��+���`a���ThI���6��VIu)�.�E:t��
-���Xs��/Zҡ�1�:��Q`*��C�c�u|���ThI���0��VG��В-����S�%Z�S��[E�BK:�<7FǷ:�L��thy��·]�BK:�<WIǷ:�L��thyΕ�o���)}��eVG�Y]�BK:�<NǷ:�L��thy.��out�
-���D���2Zҡ幕:���e*��C�sDu|���ThI�����VG��В-�������ThI�����VG��В-ϡ��.S�%Z���[�ъJ�ut���eNG��В-����.S�%Z�1��[]�BK:�\+AǷ:�L��th�惎out�
-��r�
���2Zҡ�*��:�L��th����out�
-��rM���2Zҡ��.:���e*��C�5jt|�4�Li*��.�:����2Zҡ�A:���e*��C˵�t|���ThI��k8��VG��В-ע��.S�%Z����۠��ThI��k���VG��В-�8��.S�%Z�զ�[]�BK:�\sNǷ:�L��th�v��o��|(����eAG�]�BK:�\�PǷ:�L��th�&��out�
-��rmI���2Zҡ��*��ut�
-��r�O���2Zҡ嚥:���e*��F��TtWo��gCU��'�guo�}��*Z�K�0���P�v���j�+�,��^ie���J+��WZY�n���B=�V*H���P�ymԁ��K���5��ߥ�Uך�D���k�`bxi�еf0Ql1Q��~�Z3�(^Z�r�L/���&��V\\k�K��mu1Q��z೙�	C�M�Q�w�/j����������-5�{5IV0,g�$+g����C]5>��d��*�\�vQuCA�l���K���~I�r�/IV0~9�f����2IV�&�$+gsL���)&����u���D���^�L����9��TE�:�5����U}VRX���۹�Y&����[�uȋ6�:b�TQIgTW�k]�4�Lh	R��e���׍��g}\V�~�ꮪ��yl�γ$Y9�B��-��?D+m�5�ʬ(���{_U�?ϒd��=
m���g��m��U!3�������%�K����ڵ68Wd���/�dM�w5>8OU�Q��ΦX9��R�`��e���2�������������{*//~���w���u<xsu���v������K�����å�ܥ�u���5p�s�6Ztn#�}INd/�'*ތd������P>����ݚ��bmj�Ź�$�r1]&*(����%(��1��!A9��W�t��7>��� ג�j�jaV���r�����^}��ыH� ɮ~������^���	O�e���Ӌ��$^!>�}����+���۞^t�KQ�Z�/{�g��<a��'�xދ����.����x�j�^�|�,��T�zIZ�J�����F=E�+�����>��ʓ	?���6x��x�����7ݱ7��G���������ҷ� ��r ���9 A��\N ~���@��G�����#��s�2���.D
�8���#�w��7N���$��|1��?�ȉ �O���z�W��?�}����n��s�~C��F��>�� ��Mz;h���o��O��hA�JPP �=
o�N=����mzb"Z�D���� �\�/$�\Xⲗ�������p� |�P >�( _�1�)��/���PO�t��B:� pG��;"��<#%"_ �@ ��|(�0"�B�u#0�H8>BU�	��|�% �3�H�W^Ґ9�e�d<	�-�^z�{�7ۂy��C\�>�#]�(��W0��a��0�'�W7���]��/�?�~;��mv��������?y��F�VlSU�bf��*��0�TY!�؄KZ)�&�XCH!6aƒB
�	3��R�M�����Bl%A�bf_RD����>�� 	Tn�쫢H9 9� ITn���H9 y� �Tn��� J9 �� �Tn��+J9 ���܆��B�r ���) �Z@>��0�r�R@>��|*�a�%��|j�Tn��KZJ9 ���܆�ՔJI@>u�|*�9 �Tn#r $> �:@>�ۈ�|*�9 �Tn#r ��F� �S���ȧrf��Tnc��#� �SϹ��+�X����K4���&�X~�E�Ѐ���Wnc��>�k��c�7)��b�^r������6x)_��@.4[Ѹڛ�bI��d �9I͢�V�7)Ś�f#�E{�R�0�Mi��I)��,��+I8 �9 R���P� �����6x�;  ��s��8�Ψhd�l2�,s���MX�Y�,���VK���2�"{�#0��$~��fK!
��G`>���F������|Q���7[j^x�X>�ž	����׋�#0_�C��7[2^x�X>��lux�=���|�3��
�8{�a��g6�U�q� ������Z�;г��ǋ%$4!E��B�2�C-D�D���&��h����Є<��C�"���E�}�V%`BB�n���LHhB���!Z��		M�C��>D+0!�	y ڇh�&$4!Oa@��F�0!�	y�ڇh�&$4!OA������S,Z�X�N����}��)`BB�t#��:LHhB�*��!Z��		M�Ӽ�>D�0!�	y�ڇh�&$4!O�C��S���&䩁�!h�&$4!OkD��S���&�)�h�u
��Є<��C��.��.�Nqh���:LHhB�Ƌ�!Z��		M�S��>D�0!�	y�4ڇh�&$4!O�F��S���&�i�h�u
��Є<��C��)`BB�����u
�p^#z6��z -[<Z��	'(q�1Q�V1�b���&<\z�C�<�D���h3-�/�d���N�V��hQ�ѢLHhB�C��!ZԀ		M�5T�>D�0!�	��ڇhQ&$4!׮�0�E��Є\w�C������}�V1`BBrE#�ѲLHhB.���!Z��		Mȵ��>�O��ϱG|	h�2]�I~�h�2'�H?�b�-[Z��		M����>D�0!�	�6ڇh�&$4!�u�0G�0!�	�&ڇh�&$4!��C�-[��t�p庞�ڊk�;?�e���Y���뚞���ܑ*�kE'��UF]y������g�HW?� �6���)���tkH#t���Z�:�kH�p�@�Z�@�$�<�F����A��=_"l�i���Zk@��e��8�l���+��DAS��-,fo�F�x��wZk�D�M�m򌪼�|Q����UmM]�[jN�F������C�t��g(i��#Y��;�A)0wd�J`�%��$sGzrW��#=���d�D�t��4��h��'zri�x$�rs��#�-�:ܒ�yt/��4{G��{������MU���Y3���]�g%�u�x��v�T�N:�T�.�:�E�U��鉇V��Ψ�|׺�iLy��H9�����u�|���J_�U�������C�S�O:������e���x|[dM�2+ʡm��W��O�?��S�m���g���&�]2S�ϻ:^����t���'Z�µ68Wd�����ɚ��2j|p�������'������{�\^<w�mv��h�����������/8�r��d�	�=N4���"܁�Vl��v|a2&❉�&ޝx����|�m����|��#,a��GX>���S�C�����?��Q�O���O����HI'�<��H	ܡ���	Qz�ň���M��8�ĝ��IS7ޢ׿��p����^�ؚ_�?��W-�'z�!�0ϯ�	�&���+R����1��� E�(�\I/Gԁ����M��r��r$�n���"g~9Az9"y�����$
Y�΁�_]���$��y�́H�m�$�%�LGH�^/���\�[H茐��Б��~����@�~�>��$��������}�]����n�k�Nb�_��{��w7&���&?��6��&���7��&�o���|Sx��ʇM�|S����m�GB�#����a[1?�������C�'����E6��n7�Ww�Q]����m��/��~ڻCw���ÿQ���G�ۜ��1��}�������n{�����Q�������C?:�n���a�rS�ȿ��ˋ������o�9����U�����ݧ۟�|�h���P_��q�]�����Us�?�m����ն�.���ě�c}s?���~�oO���ɶ�����D��R�vW���Gm[������e���ɀ�G]ب��7.+B0Y�M��&޹�q�/E(��_�����7�����(��۫x��=�������j�^�7���4ŻpY��(�V��/E��%x��!���n�Z:�,��ʧ�X�����KG���Z8��):.3������[���bKQ��}�P��t�_:�.1s�Æ��^���]x�0��fw�q��.<n�݅���~C�?�vv����_���>���31]K�Շ���Bȫ� ]}�\o����|���3\��+�piM�{��2mQ�jSt�B��:j���cFjmQ��]��Ӵ���4%mq F���я�E��i�ڱ{���UUp��_=�`0�ކ𰃋)�ᢽ~dQI_AL��������7������^�sSQn����˪�i�y���l���&�eVd��0;5M���v���A�%�gO�1
be�9�r���<����/�V��ϖ���+t�식��NqY<n/v����?n�d�n�ǟ6��M[�]�m�ӆ������E��1?���q��C�����2�"_����������ӱ'��5\R���*&�G?��Ji��QL�m��'��!ӗԵ������(%{�ǜ�� ���(����Q/p����)���^F�����emuָ�@�2��b�gy0ŬiN���.�2�Ch���d˯$������o~���աb��PyLt*e;�55�m|��{=du]Ʈ�`\oz�;���)�b��P������k�)�������K[ֺ�geQ�1�Ա_�{�}E���l;��'}�O�7���Ҏ]���I����(�ˇ?��z�DI4���#�wE��^yl�-�+�����	_G^�.���,�(�|WY��&�����x�f�M�Ȏ��|����<wz{�E=8��ˇ܇&����������������B��w�0/�u��Y>��<luBOy얔E���Ÿ��Ȝ�=�ؔ4U5ku���$��=�+�b\�/��m���h��ʇ#�m��[)~�{Ӎ�����[l�O����_d�w�*>��n��w��D]T��O���>�U^��]�����؟N�C���S�}���m����׫����7���$|�����ǋ�/�%
�蛏�c����wW7��M�
5�o�#����F����H�h�_�h?�^�쾫w�F�_>~�x��t�<|�>������������h�ex�ц��<�[l���4|�nt��>��w�ᗏ�ĸ�g���軯;Ǝ��3�X�I16�m)�(x2�^3��D���x.����&�_Q�Ԝ��W�����5苠*���d���������q���ק��5��L)7������-ᑼ[I�l8��4m��cR�Uԙ�_ \n!��N.����/ ��d����78q���g�q��g��^��^��ȫwK��?�5.�H1\,:ЫRz����h���'���sy�`I���,��R �e!����q��0&e�n��%�K���pq��b�šs�}U�����{U_�-op��'��%�/�ý�_�D����ר��G����.�ܫ��'�5�+�l��N�9�z����B���|p����}�n����e[�p9�>}��N�p	�|�_.yR�`�dAU�L�+1�|����)T_��u�kBe?��\�L�Z�C�W��Ն�x��j�i�0��`:�LM�
yZ ��U� ��Tԝ�;_%;ǉ�sE�:�Y�Ρ_q{��P�-#^�"ƹ$�oo�*�7�`���Ūz�������|��?x���S�����ݖ>|�y�����V|IߓV��o�ೂ�S8���S=�����:ޡ�������J�����3�wmg��G�J��	*cm���V�I��+PuF��RQ��RFN�m���K�m6`�1x�e����9J���S���nsy{|i�
ƷG��<� n�>Z���׭�Ityd���gh\]_�y�S��W�5/�c�n�����O��}}�����?�1��\��?PK
   U�mV�0��)  ��                  cirkitFile.jsonPK      =   *    