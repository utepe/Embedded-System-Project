PK   O�tV0�|�3  b    cirkitFile.json����Ƒ�_eЋ=��ٌ��d��ma��-��y���nu���:At/s�t���*�X����z�����n2�F#3�G�w�_��M{{�o����_��\�#wy�m}�}_��U]^|���<�n�|W���ݏ����}���u���2E�ں3E�V��Z7ES�M1h��>��7j�.�}�����-Am�����6�����6�����6�����6�����6%��+Am<��+Am*6W�ڄ(�c����w�]}u�K6n�뻫�������	|w��ާ�����M��jgu��b�-,���{%)�m�ȷd7��/@ �M�7��7�{�L�"�Ѩ>��s߈�x��`�����-"R�[��H�oC�""�a���v�-"Rp�7�EĮ&����R;¦ t��n���|��)���-"R�����d6���z5���ED
��dh��dh����*d_\��o�"b��o�""�I`���&�-"R c�M��7	l��ߝf��|��)��i��H��N�ED
��d����p�a�A��w-��ED
��G��P��}��"��V����]�����,t8����5mpG�,` �r^��V��O*��̷�7Y��d�E���5�Õ�U��Ec0���M��7�l���ԲED
~S��6���ED
��C���H1?�o���&�gמ����ٱfҜׯ���o��Y'N����,p�׷�7���~�s�~n�?$f���v�-"R��i��H�o��"Ԧ��l��ֲED
�p�L���^�������}�"I��"�OF'���DE��N`�/�����t1f��Ncu�#,����VwP:�����;�����t���՝��JGX�س����JGX:��X�y��t��S�
��
�;(a���Rt��VwP�ٺ{޲���Y���<H��G`����?tl�N���t� RD3>��J��c_/m� ��`�̗6v��s�|�K[R���:X>��4`���,���6 ���!���|iX��G`���
�?p��#0_�4��/X>��n`���,���F=����+��p�����X>�͑`���,��҂^�������|iG)X���G`>5�ʊ��ߌ�3�5Y(�Á��L���_�|�꬘��hp��#0_�^��~�|�K;���G?X>�=�`���,���nz�����+��яG?�`�̗2���~�|�K���G?X>�`���,��R��������|)SX���G`��c�?�?�|�KN���X>:��Q��=��9�0ͬ�V=8t��qFj,w���R�������|)�X��5��5��ǂ#�|�|t��l���ik�A�MX>��?`���&,��R�"���A���|)�X�	�G`��-
�?��|�Ky���MX>�DY`��#,��R�-�������|)UX���G`>5˕���ߌ����1��~p�������97��>�`�̗����}�|�Ki����>X>�|X�����G`��:�?p��#0_Jz�8����	��9���/צ����\Y|�axu&E^~ۉ_a�D㭸Y{'��V��V��4s���Ӕ�+�Os�,>Mr��#�~�̯tv`�����tvH�����-֖g��Hѵ��G�gJ�u�
��+��K�����9��f>�X�7\��ޞ��Ύ�\ ��O���x�z|�}�a=��w����\[~��l78ݔ��+��mQ�v(B[S��-5G��YřO_n���/7ٙ�x���B
��ۥO0�p4�ӗ��̓̈́��5EL#p0# ������Ǭ���Ǭ�˽Ǭ���K�)RB-p�PB-p�LB-p�HB-p�D��;����9Ȫ�]��LfB_TT�$l���3G:Yŏt|U�ҷE茋]�X2��+��kM�4�:��)�����l�[�>V���)�뇢�B��te�VyzV�姓�6�*�}�!o}�8�
_m��6�yzV�#�w��z�vMe��шj\�ꡳeW�79V�YřO_�z�jg�/ڡ��ݍ��B��Xg,���p>��2|Vq&�rv��*~l��"�y(jr�zj��w����Yŏ}��!"�U���u��oM���7ݱO&���ӣ�ۺ�]��&����!������WG��U|��M5��*��Tu4�ઢ��Pt�T�����泊/?ݑ/��VQ���.��eQE
�����泊�O�i,�y�ݴ�׷w�~�4����_���s�-���!	R�W`�@�Tr?"� ��1H�JQ�$H�HC�R��!	R)�����2FA�q��C��6T��4�E���mCY�}�d��m������&��FIRc$b�yo��o�$5NՂ�`�`.%I�S� &�'��%�$5�]�:�0?�a�o�$5�r��`~\��8J���AL0?���/9k�L0?�a~%i�s�h����a~\��8J����q�70?���rup#)���70?����4`~���8JR�'c��q돣$��w0&�������;�	����Q��EK�����q;z�aP:tL&ܘ��}��t�a2�����q��q�(F�0?na~%)��1�����q����6���n;>N�j������{�k�	����}˺�e�d��q��}���L&����}[]�a`29Lk��R��;�w0?���r ��`~���8JRګ�0����GIJ{�aL��[�z��߃������Vg��L�%`jk�4!�DXI�Um�i�R�z�`%V��f��K�U��DXc�%��i�9�$XI�5��D�:M(�р+���>��^���0�`%V�����K�U��DX�f�V.�W	VaU�i�9�T�^%X� + .�1�ҡ(��Z��Mk�et+u	�]2q�^$y�E�Ц��2����DhI�6���ѭL&BK2�i�ne�0Z��M{dt+��Вmڋ!�[�hL��dhӞ��Dd"�$C�����V&*�%ڴ�GfbA&.�%ڴWIF�2q�-�Ц=W2�����˴L\�e�2Z��M{�dt+��Вm��'�[��L��dhӞD���e"�$C��V��V&.;@�c�M{Det+����aZ�����˴L\&BK2�iϮ��$��L��dh��c���e"�$C��P��V&.�%ڴ\F�B���+��eF&.32q�-�Ц��2����DhI�6��ѭL\&BK2�)W��ne�2Z��M9dt+��Вm�]!�[��L��dhS�Z��L��dh�޹GH���e"��ß@c5V&.�2q�Z��m��"�[��L��dhS��
�$�J&�Y��lzrJ	2q�AZ����ˬL\&BK2�)���ne�2Z��M9�dt+��Вm�E%�[��L��dhSN-�:��L��dhSn0���e"�$C�r���V&.�%ڔ�MF�2q�-�Ц�s2����DhI�6�ΓѭP��9-b�F�V�j�ԭL\&B;?��:�����e"�$C�r2��V&.�%ڔ[RF�2q�-�Ц�"�-e�2Z��M�>et+��Вm�Y*�[��L���h?����ꮳ�B[X2}Q�:�W��N�o�.�üR�BnڕR�ɮ����{�{��R�;ܗ[)e!��J)��WJY� �R�B��V2^��.��V�~��V]+f�Ԏ�b0&�t��Z1#ޞ�9?�e��{���q&k�lO����V�h��׊�x~6�Z1+^:r��ъ�r��d��s4֊�x~��Z1O�xzZ��V㋗N�(�m\��,(�]a}m�ʶCښ���n�9ݫɒ�a9�,dI9�*x��:4��W�m(�Dm���l5�|��r$K
��eI�2?�k�s�gI��,�]�R�ɦ2K�ɖ2K�Ɇ2K���^�թS�7O��yb�)�'Ɯ�ybF��V��xŪ�]��Lt�&�EE�K��(��Μ��YRN{__ծ�m:�b��IT۵�kUe�9RN��ee�����Q��v����!��M�i�,)'YHyt+8����hU�����{��O�dI9]G��V}�P��ꦨMp���Ζ]_/�^��`XN��޴��vh|ԋQE��]A�u�R�:
��(K��7ʒ�y����!4ʫ�9�r���鄢&�>졧6~R�u���%%�387��eUE)>�V]���[ӻ.z�������d�����ا�mr������0��t���:͒%�$KS��ʺ0U��ઢ��Pt�T���>�����dq�ˮ�UA�G)����}YT��Bt��Ω�,)�,?�b6�������x��G���J|7���]}�˷�$-���@�@��� D Aj�e"� 5�"� 5�2"� 5�E"� 5�X"� 5�k"� 5�~"� ��#1.�qn�	�Q��6\�0�|7��7J���&��&�GIR�	%̇̉�$��T�	��5̏�$��$�	���u�a~\��8J���5b�`~\��8J��΂b�`~\��8J����b�`~\��8J���c�q�70?���r.p#)���70?���r���`~���8JR��c��q��(I)��	��-̏�$�\S0&��0?���r��pc�Aq��0?���r���`~���8JR�yc��q��(I)�l���̏�$��0&�w0?���r��p����M�w0?����zØ`~���8JR�[c�����Q��^V̏�0?�$i���پg����Q�Ta%V���yFK�U��DX�f��-�W	VaU�Y*�T�^%XI�5�]"z����h@��DXc?HD���SH��k죈�u�v
�	VaU�Y�)�T�^%XI�Umf���R�z�`%V���BK�U��DXӚ`��@&��%ڴ�YF�BQ�P�%w�L�E2��-�Ц��2����DhI�6���ѭL&BK2�i�ne�0Z��M{dt+��Вmڋ!�[�hL��dhӞ��Dd"�$C�����V&*�%ڴ�GfbA&.�%ڴWIF�2q�-�Ц=W2�����˴L\�e�2Z��M{�dt+��Вm��'�[��L��dhӞD���e"�$C��V��V&.�%ڴGTF�2q�-�Ц��2����DhI�6�ٕY�$��Вm�{,�[��L��dh�j���e"�$C�����Vh���rE�����eF&.�%ڴ7_F�2q�-�Ц2����DhI�6�J�ѭL\&BK2�)烌ne�2Z��M�+dt+��Вm��!�[+��Вm�%"�[��L��dhSN���e"�$C�r���V&.�%ڔ�FF�B;Ʉ����eV&.�2q�-�Ц�A2����DhI�6�>�ѭL\&BK2�)���ne�2Z��M��dt+��Вmʩ%�['��Вm�&�[��L��dhS�3���e"�$C�r���V&.�%ڔsNF�2q�-�Ц�y2���!��C&.s2q����DhI�6�2�ѭL\&BK2�)'��ne�2Z��M�%et+��Вmʑ)��R&.�%ڔ�SF�2q�-�Ц��2����Dh)���Q�]��:[!��%�u��|e������9�+�,�])e!��J)y�WJYȼ�R�B��R�[�����z����+�,�|^ku ��X�ҡ�k�`�w�hյb0�t��Z1^:&t��k�/���VƊ�N�\+c�KgA����׊�X�ҹ�k[]�/��QL۸��,(�]a}m�ʶCښ���n�9ݫɒ�a9�AeI9�=y��:4��W�m(�Dm���l5�<��,)'��%�^��`�r��dI9�e���t2YRN��,)']L���&��@Ƌ��ӽ�<1�=���s҂�
�u�.��D�mB_TT������i/�%���U�J��3.6(Q@��tAu�]k��QUFK�#�$KYV�n�-L5kkg������b���ԝfɒr����AW���QJ��QU�jh���!��4K���u�Zo����n��W�z�l����2�%K
���gmZ��E;4>�Ũ�i����:c)T��v6G�iO�#�F'���U��U9�E�tBQ�K��S?�κ�zɒ���B|����_��z]���]�K�e|�YRN��O��]���69��EOc�P�fh:jz�^�fɒr�����Ve]���_@pUQ�a(:k*��l�QGYRN�8�eW٪ ꣔��Eо,�h!:]_��Q��]��.���{{}{����v�N����Ww����usu�������w_͉�X݂o.Ϯx=ֳ=�s�zv��_���X��ю7	2�d{5��h{$��B�hF�j�5#9�\u�Ʃ�8�r�]fF�,%L��pP��1ݙ�AٳӳN�ƙ�+?~}S�kI�:i���B;���}ɫxGܷ�$z� ��/v�r�~���1��-���x����������}��<>�o_�񬺯X��jqRJ�w�|:��1]��<�ǳ���/|t�=g���9Q3�����_-��(&
ACT�q�X�Qf� GV�1�1��<.�Bt�br�,Y,��7,�Ф�߾%�_3��*&sV����A%b�3W�8�������21���4N.��0A�2K� 	��<�X/!��"`��1#��I�ϸ��TP��O��q=�q��~�<C{�w�׾��7ݡ�گ#h�����8e@��\�� �<6 �9��' �j�2�|r� Ч5�=~:����>]u!\0xq��W_#0���BTw��Q�WY��'B/f��4,{��g̬p�?����è��6�B�j#{���M��Z����/���	1�.^a�U�B�����x;v�{]O�����`��c=���R/�Z�S�{���XL� ��P ��( +�0��]h����P_*w�����P#lT�pW"~�H���u� ��_�ȇ �R蜷X1�,��g��O`#`8���̉X�U�x���g����zS̗�]v�� �>}e��)�O`-*�À^�z�ҏO`�h+����hm��:V>z9+`%����=K�q�s�ʃ�'�Ϳ-��0/��C�]H�d������Znr:��=6��:���#x}�"�n��! ���*�"}�J����"�y�����?��Ż��o�a�������x�#�y)�܆��-b���I���<�L
�5�dR�E�14��-B����lj�Gͤ`�Pc>k&[��a3)�"ԘO[��㮜 '�fT����Ţ9V��8�1}��3� ޗ �/Cm�s9 � .�/Cm���r �0�0_�ڞ��� xbb;N�P�3���7��Հ�,_�ڞb�� �S�|j{���Oǃ���=�ZH[�\,�{��Pۓ�&��
mEr��9k'mEr� Η/Cm���Ƭ �k Η/#r �/_F�@�% ��8_������eD���ˈ��,_F� tf�2"���e�������mEr� �/c\�4�C1G4,��Z3�b��X�H���]��L��|1_�8E��[�k� �̗9 ��/#r \3_��8@W�/c�\83[��#mEr��f��q ���ff�� ���]�bms��H.ց1
f�{@${'$�͗9 ��/#r <5_F� xj��)��/#r z�|�0(1���1s���`3GVr�϶�`�g)��jCSzf]��%��|��K�џ��G`>�1`����|�QX�?,��b��?����|��_	����|j����`�a�̧6XXX>���1����|��@������E������� c		M����uJ�Q	:,��J�
��pF8���;���i0Z��XLHh´��Ct�&$4aZ��!:f�0�G���		M�ֽ�u��]���&Lk��:D�/`BB��h�c0!�	�^	�06:l�P�ҿ@bt�[��j��*�C��
:N��8E��0!�	�� ��q
��Єi_Z��8LHh´	�Ct�&$4�����
��pF8
c�P���?���0�<����gh �ht&$4a�t�^L��b���&L&�:DG1`BB�͞h��0!�	�FU��+��K��Q�AG1ŀ		M�6�u��b���&L���:DG1`BB���h��0!�	Ӧr��a��ЄiC<Z��8LHh´��C��S���&T{�`t��S���3}f[�X+�����J�a˜p�fNk0pJ �V):��p��h��{\��\�Q�EG1�c�����b愓[�
)KZ��LHh��CtP&$4aJǂ�!:��0��A�Ԁ		M����u��A��Є)�Z��LHho�Ct&$4aJ���!:l�0erB���		M�fǧBbt8#�D����j�]�J�a�p~t�S�(ơ�0!�	S�2��Q��Є)�Z��(LHh"��ŀ		M��ۡu��b���&L���:DG1`B:E����Y�ƕ�g�מ��,?�%����ߚ!�@�ׅC���͒��,?K����,����d�k��m�\�����V �B�gѭ0���V ��Ƕ��5D��{����ۚ�3���~�!��O�\���+��|�\���F=?�k�������[�ea�K��/@qZ���Skq�m�����Pv���-*�Ehk�Bo�9�u�*�}���!�����{=ԡ�E�*lC�&�Ӈn�d�AW���q�EX�Y�g��в���ϒ��w�۷�qe�;u4�JqG�۬�G�۬�GZ۬�G�}y�x��|s���ͱ�'0/��<ys�^��y����8��A�PV�N�`��7�/**]
b�yݙc�;��1��ڕ�-Bg\lzb����`��tM���-GN�#�/��֍���*m�L\?uB�]�c��*���������[_4���WC�����Ǟ�U���]����2�[��	�P��ٲ���������i��i�3������FM�w5�K��(��*�?�<��H�c��*~z��"�|(jr�#zj��Yw�����~�B�.�*���%��Eߚ�u��o���OV�#Ϗ�o�.��z��a�'0C(L345=y��=?����7�ڪ�S��~����C�YS�Fwd����*���|�U�*��X�5u�/�*ZR�������U~���./>���6��(���ݏ9�Ż�/R#���X�)u�RC���R_8u`S�s�+�=�qtol��)�1��7ḅ:��c�S�1�թ�N%t*�S	�J�TB�:�0�Dj��������ǂ9�1���rۏ�K/��:��i��
�?�H_eI�^�`帷��N���9d�@��W ��)?����y�?��s/F1���h�����D&3s�	�����ڽ=��LN�����kw@�����2����(���6�.���!�밢n��blW篣����Y�xsG_�㸯Ê������X��k���o����L��fD\oc9��1g:`�D�2�Nw��+�s�X���w$�u�9�'��&�P���� N5���W���x�;��d�:�9�g��9���H��F�������<���gj���J��n�D33L�H�	K.!�ܜi2�y/���.x���?�{�\�M��}��_��x����%�t��/��Kf~I=]R�K�t����%=��.�����R5��.��%z&�9"� `�O����3>���YW4W=���:���с�=�8�ߜ�ߜ毮�_]x�g=�\��l%47����C����z�c�W7������aSʱ��l��w��&��6������%��u?<�a��̗���W�C�����/�n?�wW�8��݇����%GE�?�]ݤA�����{�zy����1�����2����*�_ğ����_F���������?]�_5�������|��뻋w�=bE|W�<u��x��ؽm��{����D��!��n��.|U��vG��eT���L����.��g�)�s��V�E�b�U�����1Ҽ���o�m��9�ˋۻ�X]����C�S{u�^�O�uQ)��]�*Eؠw~���.xx�P�v��Y*AK%�B���_�^.8�p�.��K%h��%����R�/�����^��+j犯���>_�p�-��K%�R����.���}�/�j��¬�/�j��¬�/�j��¼҅�?u�[v��n��������w�����������/.�_\u�_�
)WMla��U��4��T�m�x��׷�a���w׿y*۵����FU��m��T(��ZG���˦���m�����
|���d��;���s�\�R�77v
�un膢7i�m���tA:�kck��/x���?�I��N�?���o��o�����6���^5}�Q�u]4&m�z�u�=U�����}��C�#%�J��i�C�����b���:�; �׷��.�ҽ��RA��Jj���jW#cS=�0<��������T.����z��?Km����܌ǻw����,�<�����/vo�����]w���?	��.�v���u����B���6V��j��W��^=ֶUu�}O��ՒqFWC�_��,l]Ų�nm�aZ���!㪣\�+U4��T}\�c��hr֨R5��EN�U+���X�5eQuu�8:m�n�.��q�j�������U��x����Ǜ߿�y�����M|ܛn�Wޤ��|����on��=޼���ۻxw�����]����]}us@�]�������]a[���}�e���R]^l=�oS���Ѧ�&o�Zп\=|���]������6���ުh$�>�W��}AΕ��}������7�n��ݎ*�d�|Y��6*�ʽ��&~5]�K�����f�:v{���M��ӾQւ�iߨ���f�;�լ��6Ho� ���e�|�<7[��e��6��ePO7����^e���J��F�̨�O��~ۖ�ǫ�7���S��nk&���nS�z��/C�^�Z�TGz�䂮��5CѸ�*�@:�_*6�uS�.�����\�R���x���OX�dITƞya+��j�j�/?��������z�&�|Ӌ�>]p;7M�u�>_��_.�i���M��4
x�u7�\(�_������xA�������������t>�����:x�lI��b��K
�ڿ���~(��[�b��b�-c�oT_Qזzq��P�a�ĭ6��eDK�ԎF趿�<V��ϼ+����_�������y�l�̞MT1f��)tcCQ;u]�F{P�wM�����Dֲ���a�G�dێ;;�"n*��/c���O�H��o��&R��Z�a��2�{UE��詥ٵ��V]l{}��!Ν���M���2�?���,{���M�!|췕a�scط��<|��*�@�ӻ���ٗ�����Ƙ]����_}�����?���e�os�ã����å�z�O�����K��2v�*�[bW$� ��q��}t6M3���n6�/����&s�Ǒ�C��_MY�T��{��C�}۝��nS-����M/�Q^*����I���0��K^u�o���3�������>v�ɻ?�^�wS���?�|�룱�M��!U��8�V�Roi����g��g����4�q�g����k��7_o>�o���|�{_(�.��t�e����^��'��d�Ӣ�4�YצP6ڴs�Kݱ�Z�V�������:ǰ��a;�۟�i�� �[z�lc�Z��c�c�;�A���)$��SM���/��1�v��+�_�m��i���P����.b����t;����շ3��6�l�w9k]����Ӆ�;��Nl;´���r:��.k����%3��z�o��ˠ��+��?��Wj�P�V�JE��1�H):j
N׾�6�e9p23߼����S?O����}7&��/���-��e4��/����v�'�ɽ��m���11�n��Ǟ�3}Z����d��2��Y�jalg��ė��]�`I*M��{33�����z()�<��AG:�픅�E���ϵs�!]!ڪ*��=�w)�^���U��m����}H������ސ�KM����Y����%��}���B�/�����t���2G��1-:���W��K��[�+=������yZ�r�V��
���(�n�Q�]��WH�(��r�n�n���e������������t᫱��O}�u��q��G;����|i��C��P��mvo�7�6:�P[��}������]�=��4;��mci�m��,�߶dc;$Gm�LG�lmb�Sv���l�����Vv�J�w��4��]U����Uof��������Y��S��w���o�3���*z�2��w�=4�6�^����6�l[�?�6���lۜՆU�ƨ�&S���u��u�m��ט���qnM�,o3�G�T���drWns����H����I�������.{��qs���� �5m.�H�\4��Y�B9���]�?��Yg�����Kf"0Qc��0�߲�u�#Ҵ?s�m����+]�hs1@ߢ�Š}�>�\LV_Ü��x�
�̤'Z�`P!*x���e�B's[~_��}�6�F�\,��\��װge�^g���`�?�
^��w��cc6������VW���}��|Z�'T�\�س̥��Lf�������we���?���ɑ���(9<N=�T�;�O���#��ͼ�O�T�{Em�D���g��fjr�+�`�� ���`�i�q�Ya瘛യ��;+�����a�E�gEc����Ί"^�z33���/6�����i/������ �����"��ۖf��2kB|���!���c���]+X�=��k�fЉx���]�;�ۻ>z�����i�MGaM�$M�D���]��܉��偻r�;#�X{��������
T���gFc�ٜ����ͼŚ���V��=��\�O�xҾ��<�ٿm�^7���#�.N�In��<����V"$�<p�E:�Tl���e�k|���獷��g0�}�"�����k��>��mit�3a?�-�BY�}�6��O��O�/�<k�s�<�S�������3n���0<-�̱�u�T���s��ژ%:�`&����;���3n���q���	����O��0�WS�f��m�Q�s�L����59��[�!��&`�܉��:�D:������7��k�e� w��z�Π�/�@�$�_�=��&`M����]��4�x��ۖ�)Q����������x�,�~��������������~���������.~��PK
   O�tV0�|�3  b                  cirkitFile.jsonPK      =   4    