PK   `�tV3��Ŵ7  �;    cirkitFile.json�}�n%7��4��.��a�Lֿv����1�Y�6��F�j$U���h_f�i�<R�N^�a���T�v͠-)����`|���������ۻ~����������ˋ�����_���۫�����/w���.���~/~|��]_w�m,�SD��;S4me
�uS4u��v>P��z�v�����^�/��Ԏ���N�1p%��ac�JP;�����v���+A�J6���Q����ooo���]W;���Cma��E��(HYo;E�%�<���b��+AE-<W�����⮾��Evoo�뻫����/L���T��Ĭ |=���=i�]��`oo�z��<�""
���Q�����?��ED\?N|,`��(���"b����"T�( Q7 �֜!1�h����(����X��f��(܁� .%s�|���.�-"����F{dp��Ç��5��q��E�?�E���El(b��(�C[DD���?$�ED�0�8��0�
c���[DD���55GZf�t�-"���p������*�Ph�����?[DD�F#��C[����6�`�V}�O�tU����e,t6��!�FI���� ,cXN�����Ǹ�?rZ���122� ��!��9s��}ՙ���l�e��(�#-[��9>[b��(�իJF�bN��;���q��]{n���c̤9��Ɗ�?�;ְN�q]s�u��Xշ�pٴ��i�g�l�f��(��4[DD��wǆn�P��?�ED|��Q�gHg"�����w�B�С;d!I��@�XH��	}2:Q�D'0q����EGXt��bu�����#,:�3X�����.�|��,VwPt�Ec/��VwPt�E#��J����N�<Vw�;(:¢S�
��
�;(:¢S�w�#t�����C����zF7p� �5��#`���	�������RD3|��J�Iɱ�K'M��S,>�Kgd���,>�K�{��S,>�K����,>�K'���S,>�Kg����,>�K����S,>�K�����`���G`|�� X`���G`|��#X����
�h0��`���G`|�'X`���G`|is0X`���G`|�,X`���G`|jv:)��>���d�-D�`�2=��V?���񱚳b.>h0��`���G`|��7x
��`�_:����`�_:f���`�_J �z�z���0�1`���G`|j�)����Õ1D�`�d��	����R�����	����R���������R���������R���,��`�_J����`����6�U̙�i�����g��3�c��ְ�K)m��',>�Ku��C��A�'&NL���h�ٞ�{PׂI��&,>�K�����&,>�KI����&,>�K����&,>�K����s`҄�G`|)�X`҄�G`|)gX`��G`|)�X`��G`|)kX`��G`|j��)�?蚏��`�����/X|���l�H�,BL}��`�_�K���`��:�f���`�ͳ�1]97�A	fN%�9a�_J\��9a�_J���9a��	|3N�nnM��+>�t���4W��<��,���2��,F����'�U�i�ٍ��� �X|�<x�0̅^ũ{`~�s>>�M���'9�'����L5�.xk�i>���7�l-��w�kq������~���Z��h^�]ع�.sf^%�ߚ]\��<���n\�~sg4����z�X���ϳ�掹���5�q8������z`�6np�)
eWX_ۢ��P���.(�[j�Ђ��̯������n#s#/��n�d@��o��3��c~}�f�/'4rgn�b�����__ ����Y��ÿ��ӫV���%4�^�%4�^�%4�^D%4�^���c}�}�T�〬
�u�.��Da&�EE�K�F�^w�H0�U|=(��֍���l�L\?uB��+c`s��Y�׿N�۠����C,���qT�ڦ�m�?����G!�z��hYTF�66cm�+T=t���X�c��*���z�M��1�h��Ǻ���
j�3�B�Q8>��:���L��1��U4wUua�65�d�COmP�ű��Yŏ4�wnrYU���5��^}kz����tǺLV���Gs�u���&��6��!������WG��U|��M5��*��Tu4�ઢ��Pt�T�����泊�ݑ/��VQ���.��eQE
Ml���泊�}0U��/L�!q�PTC��5-�.Խm�Y]N�#V�ڡ�]Y�~p�u]䜵
�T��u�Y]N���+j��i�":�2vؾ�Ί�������)u��Y�ǯ�<��=�����ۻ�7?q�������s�2��]�$H%/�A���� 	R��b���H1�@�Tb�D Ai�-
�Nn�4�G!�P:	J�����0�D`r����l6�ym�ۆ�m���0�<7�\7J�g@�`ޛ`�%I��� L0N �K0Ij\a�yqy_�IR��;(���q��(Ij\�a%5][̏�%5MU����(Ijܞ�$����	��5̏�$�ّA����q]�B_����Q�ԸD�a~���8JR��
Ä�I�M���q��(I)�'��x����	��,�K��z&&X<�����0����{_���I̏�$��@����qk��E��11���G�[V�3̏[�GI�~�8���q��(I)[̏[�GIJY�`K?0?�F��S-�8�w���w�cb��q7z߲�t�21���{��u�q�ín�޷�UX3Y�(	�;X<����t�0�����q���N�	�`�r,��a~����(I) ӊ$�Q�E�>��hg�#���#��j7Ms�i�i��T�J"X�n��.�W	�$�U�	�R�z��J"X#���4� FXIk��D�:�#�рV�c�N�b4 ��D���4k \*P�XI��M�	¥�*��D���4� \*P�Xi+��IB���b�:AK2h��f�
�.!�%ûH�x��Z@��*A�����V�}��%�iϼ�ne�Z�A�����V����%����ne��Z�A��b��V����%��L��ne�Z�A�����V����%�錏�/AK2h�Y%���2�$�6���ѭЊ�В�/�2�L��2�$�6���ѭ/AK2h�Y>���2�$�6�I�ѭ/AK2h��J�����9F�錨�nex�ZZF�_��2�L��2�$�6�ٕ٘$��DВ�t�XF�2�L-ɠMg�et+��DВ�t\F�B���+��2#�ˌ/AK2h��|������Vm�1 �[^&��dЦ\	2���e"hIm�� �[^&��dЦ�2���e"hIm��!�[+��DВZup�R�2�L���+�\���eV��-�E�`"hSn���2�$�6娑ѭ�I2��d2�����m(%Ȭ�-��[^fex�Z�A�r��V����%�)���nex�Z�A�rQ��V����%�)���n�/AK2hSn0���2�$�6�8�ѭ/AK2hS�6���2�$�6圓ѭ/AK2hS�<�
e��Y/A�n�E�V�����_k�N��9^&��dЦ��2���e"hIm�-)�[^&�����}B)��J^&��dЦ\�2���e"hIm�Y*�[^&����~�#����]g�!���d���I7e{�)�-ٵ{�7JY�M�Q�J6ٍRV�xo�b��Rܲ��(e%��F)+��7J�g���y�Qʘ�y~��V��w~=�V1���o��*c�k��n��:~���[;�����ڝ�[Ŭ�A�*f���}-[�ޣ�^g�U��ƈ�-�[�`�x�˭b0V��r~7�V1��/��*�ъ��hl3Z��ꋭb��Oo��:�b���?�i-�)
eWX_ۢ��P���.(�[jNG5YR0XNv�,)'���z�Cc�>xU؆BLԶ���V���'���#YR�Tl�%E������R�)�%�B��rw�F)'��,)'G�,)'�,)+w�l�:u��扡S�7O�>�}�ĘS�7O�h���}��9�W�
�u�.��D�mB_TT��TG�^w��͒r���ee������6�v����!�fW���4�,)'���6�**5����hU�����{��OcɒrzTr��z苆�X#���6��:[vu�^FeI�`99Bz�jg�/ڡ�Q/FM�w5�K��(��Q���5ʒ����1��*v!Uua�65�ԙ��ڠ���^���ni��b=ʪ�R|�V]���[ӻ.����YRNb�]��]��z��]����P�fh:jz�^�ƒ%�$��B[�ua�:��ઢ��Pt�T���>�������ȗ]e����RZSA������&ZA��FYRNbL�F��tH$ �P��jMK�uo��͑r�vU;t�+������ԤvC��6���2l7G�I,��&z���^����o�Ǥ8(uU$U��,YR�c�y�{���?��ś�>��~�X�wӿ{������~�Hо�B��q�� 	R�xA�F^A�F�A�F�A�F�	A�FA�FNA����"q^�a~�`�%I�0�`��`�%I�'80�`��`%I��0�`>�`N%I� 1�`~\��8J��/Nb0��o\ ����Q��~�	��5̏�$���0̏k�GIR�uk&��0?����+�:����Q�R.J&�L
n*��̏�$���0L0?n`~%)娃a��q��(I)'̏[�GIJ9�`�`~���8JR��Ä��M������q�����	��-̏�$�\00L0?na~%)��-������q�����	��̏�$��
0L��M��&̏;�GIJg�a�`~���8JR:s���%̏�$�3�0L0?^�������ug���R��jRI+�`U��Yp�T�^%��V���GK�U+�`U�Yn.�T�^%���ȻD�:K�рV�� ��RrA4 ��D��ED��t\H`%�j7�Ņ�
ԫV��v�<\h�@�J`%�j7����
ԫV�����%��dЦ��2�b]B�K�w��"�%��dЦ��2��a_"hIm�3/�[&��dЦ��2��aa"hIm:� �[&&��dЦ�2��ac"hIm:S"�[F&��dЦ�12��ae"hIm:�#�� ��DВ�tVIF�2�L-ɠMg�dt+�"&�$&�˴/�2�L-ɠMg�dt+��DВ�t�OF�2�L-ɠMget+��DВ�t�RF�2�L-ɠMgDet+��DВ�t�UF�2�L-ɠMgve6&��2�$�6�=�ѭ/AK2h�j���2�$�6��ѭ�nE��2����2#��DВ�t6_F�2�L-ɠM9dt+��DВڔ+AF�2�L-ɠM9dt+��DВڔ�BF�2�L-ɠM98Dtkex�Z�A�r���V����%�)'��nex�Z�A�r���V����%�)G��n�N�	%��eV��Y^&��dЦ�A2���e"hIm�}$�[^&��dЦN2���e"hIm�E%�[^&��dЦ�Z"�u2�L-ɠM��dt+��DВڔ�LF�2�L-ɠM��dt+��DВڔsNF�2�L-ɠM��dt+��C(͇/s2����2�$�6�2�ѭ/AK2hSNF���2�$�6喔ѭ/AK2hS�Lݖ2�L-ɠM�>et+��DВڔ�TF�2�L-��pUtW;���Cma��E�k�.���S�[�k�0o����v���l������(e%��F)+��7JY�n�Q�J>�RV2Ho����y�Ձ�c�k��n��ߵ�U���X���[�`lx�Эb0V�1V�v�V1+^��r�����UƊ�n\�*c�k�nu1V�v{�1m�����Pv���-*�Ehk�R���tT�%��d�ʒr�?y��:4��W�m(�Dm���l5�<��,)'��%�^��`�r��dI9�e���t2YRN��,)']L���&��@Ƌ����^�������Ĝ�`��w]��f0�u���.1�Q�ם9�e���l���l�[�>������CQw!D���8��ƒ%�$R�]E�����������6}oC��i,YRN�J��V}�PkduS�&�B�Cgˮ���h�,),���i�3���������댥Pu2ƶ)��C�L�N��!4ʫ؅T9ԅ��P��Rgzj��κ�zɒr���sC��(�*J�Zu��oM�أ�.�7fI9�%v![w1��mrv�k��Ba�����{uK���X�jmUօ�������C�YS�Fwd��6ʒr�#_v��
�>JiM]�ˢ���huNeI9�e0U=�/L�!��PTC��5-�.Խm3l7G�i�U����,Z?�º.R���w��뺯��͑r����ޡ+��,�g���1)J]�@U9�2�dIy�������b%n�o�vW��.����⇫��~�����iwu�������7_�᛬p��KƷ+^�������o�����m�bT�O;���d��Ő��;@®JG3d/�Z3$g�7��qj!��\u���",%L��p�0�czb���NϺ�g/���Cn$9�z�W�+��G�}�kxG��G	QDn ī�j���>�s�d�����[����N��������|>�?o_�󬶯X��qR�^�c~���.��\��Y��W:]f�,i�Ú�u��1����PJQ-�-S`��Fά09�1$gy\���,��岰L%�TC���Mȿf�W�4L��+K�\8P�	嘹�����¶ݖ��u���r�L�n?eM�0C��,�v	��"0�4;�<\q;��TP�.��"ͥ8l[�N��<�͚LׅRF���*vsp�Μf��9n?���<g��yV��S�1�=ö�3ᜏ��xB�YK<�	��	�SqPUm?R��<sV<��g2�i����v����ۿ�ݮ�閶>}�Ǘ������� ��� ��� ��� �{���[�^�|���Ok����i�G����;� ����i+�< D�q�E�"[���;�� ׽�vglS[p�	[��0C���7�Xkd�/��G�� v�r��Vw�0u�[Z���5�K�Q 6�2ǎ�����e�6"�⦇@`퇄����V8��ޒΏ�;�( �( ��( ��1��ݵ���P=��������"l��n���H���M� ���������9o�?�1 ��3�
�'p 0������	.�"& j�D��>/rxӳ�g8�S�/(kI�8���;����	esO�m�9�G�>؉ }���y8	�s�����Ij��_�s�Ǒ0���� �L��I]��(�-Ng���V4^f�c#�G/�VD�����ě@����9�1��s|�	A��N@�v��r�M�Gj��;a�p��'Ɓ0O|B���'�/�!����'�"[�^�.!���(-�x��P̣�g����biT���S�.�W�ƶ�A�l[��l I���(�9�w�u������?��ś�����s���ݻ����Ow������������-B�w1Q�E���$&
�5�'�D�����(�"�x�![��CT����|P_5lj���P5�3R��Լ�Xg�h/��k�v�~r�τ�p�|j&���e����\ /Ll�I j<���S@���A�� �U�+_�J3X|s���5���2&��j�m�2ƥ�i��,�Era�/_Ƹ<�X��ɅU�a1'/4�5k�k�ˈ����2"�k�ˈ8 ��/#�@�4 B]p�|*M[�q��f�5 �˗��|*�܁�y#,@ ̗q �-_Ƹ-`�b��ڋ��8_����,�bN�Y�/��V1'�,b��#n�!��� O͗1��D���-�S�eD �̗q \3_��9@ ̗1朙�-�@�^$ւkf:p�n�53Tp�n�kr��"��f0�\xA$;A ��ˈ8 ��/#� xj���R�q,�2OX� �͗q �h���0�1��>)?��s|�4�3����.�~�H�^�h��ٖ4�˒G`|�w�^�?����π���G`|���g����#0���������#0�C��W����G`|j����`�a���U`�U`�a��z�C�� ��,g���g��36���g�?7 �"$4´��C8)��4-�殁
��p�p��"��Ӗb�J�\����vh��|����Vn�ќ����A�
�Ѽ�p���_e4u!4w#$4´��C4#$4�tt�C4�#$4�t�=���-`��F�fIB�1:D�0B5K_��!|A�S4��h4O#$4�t��C4O#$4�t
�C4O#$4�tb�C4O#$4B5K
����d*��CXd�ŨM[��Iq��<Ch��,����	E�f4�#$4�t��C4�#$4�t2�C4�#$4�t��C��0��04�1hc�,����,�"T F�3��-̋����Ih�JѤ����)n�Ѥ���ӑs��,����qy�Ѵ����Q�-����:��C4m#�_;;��@�fW��U�f1s�0/BN�!�*E�0BB#L�,�:�y��yA��&5ӻ��UF/��N�oY�"h��I!���'h�I!��d-h�I!��D3h�I!��$9`:4�#$4��C4�#$4��C4�#$4:	�C4m#$4�	�C4m#$4�
�C�i�k1�\�N��*E�0BZ@8i#�� ��84�#$4��C4�#$4BupF�hF8���x��(Ѥ�D�0BB#L���:D�0BB#L���:D�0B:�p㥤�$�[�f��%M�X~�xvc��|����Ŗq�����2�n,?�F�n�>~����ݏ_������0m��5���{[� o0K*�U ׄ�w�m0K�U���*�˛��a�����f{x/�Vy\��߉�U �l�;��e���{8�a��/�2���VG��&�8�u~��VG⌶q��MYP(�����m�"�5u!o�9�d��~�H��*�Ky��:4��W�m(�D}���l5��-���p���H�%nᢄ�%�d;�,q1�J��w�Jč��Y双�Y��Y�g��i���<y�ͱ��{��|s���u���<y�n���y�n�Xi��w]��f0����.1��C^w���*�s�ee������*�v����!rnWƁ������>)o�����|��QU�jh���!�������\����2ⷺ)j\�ꡳeW���Vy�����޴��vh|��QE��]A�u�R�:
��g�?�?�<�����*��*���]��\�COmP�Yw��Y叵�wnuYU������^}kz����tG�OV�#ߏ�o�.�K�M�(tm�GC(L345=y��}?����7�ڪ�S��~����C�YS�Fwd����*���|�U�*��X�5u�/�*ZRhb�����U���S�����R��j��B��%߅���Q��)��T;t�+������ԡvC�j�������?�}EM�pWDV��۷�Q�*�U�:�������|y��U�{��E��o~��!Po��HAL
<R���t��>MP&.��u����S���=.׏��cJ�q�n�iЩ�838ο��f�aˑt�kM:�Щ�N%L*Iݷ�Z�g?̉FP����	6>|.ȉ
��r��C$�e:���-�e���9���@�=(���
丨�Jg���9N�Y������M����.>Lb����*k�j�P�Z��ȚW�T��+O9T�5|��݂6S�5k�Qe����(nuXĘ��P�V�5�����#��:�[δ�ڜB����:�[֬�]@Tq}��y���H�vae�ʜ1f9Ok怈�m,ǞY��L�Q/sw����=�j��y��4'zb�n�o=-�A2�f�e���?���w4q��]�s���3���N/��#\���i�#�\?x*���hf��i��9��y��4O뼍����X�B��y�j�N��ȍ�q��뛃h�c7�\�Q��7p��C��O�����(nI:���<�0�6�2���Ä�C����u���i��w����S��*�!L��Gv��<>2�G��?��G4���#����U�������(��B�C��0��g~^�	>��ӓ�h�,zR1�uLO����=Վ���O���{�%͕IO�@sS�Oj�s���M7��~��^��S�Ѽ���^�\/��z^�T��C����z��'^������qZ7�[�f�w�{������&�?�'��q~�%>�����~���~�����������{����LT�����M�)���O������ߥ�~�TZ&kxws�_ğ�ዛ�F�o�����������j���������]�]�y��M�}}�n�ۇww��1 �_{��{wus@������6����W�ko���:wQ�	��c�m��Ye
�*�UmQ��pUc�_��v���o�}����ˋۻ��\��Ż��O��]{�?6��E��kw髈(���/޿~<�P�v��Y+Ak%�J��>��?p~�]+��J�J	VJT%E�9��_l����	=��=�U9���O+�Z	�VB���)��AYM���`�
Of���`�
Of���`�
�歐���K}���r�����˟���7o���������o.���/N���+���������CaB�J�T�m��~���׷�a����׿,۵����FU��m��T(��ZG����l���r����UUt�\a���<-���m�{����~���óºi����MZQ�-� ]D ����5��
����_�$�Q'�<��5��wW��3��6���^5}�Q�u]4&m�z�u�U�����}��m�LJH�Z�E�D�dM5U5t��;2�wu�� �׷��s4J��:K�>*�����]UP5hS=�0<��������T.����z��?K�����܌Ƿ�?�ӓY<z�W��O_<��ۻ��t�]�(��K���]W���a����W�ml�Ԕ�����W��mU�x�S�{�f\����D���M+�U,���6��ޙ>,W�*]�����z��B�G��F��Y5.r����x]]�®)���c��i���жǍ������_o��W��û������on^���z?����ww�'��ۯ�����W����ݼ���ۛ�v�����]��.�����Ys׿�뇾���=���}�eD�󥺼�{�?$���ѡ�&o�F���z���]wu�o���~p���ZE#��D_��
r��@T�����?>w��L;"q)�<*���q8Tƕ��&��.���|�Qt�UÞ6���j���46��w4����n�ё�fa�|���������4l��c|����d�����qܫ�}���Z��rߊ�U�	�o��r������o�w�L�5��!�U����2T�֌�걍�s�����E�����8~�8��M]�/�O�\֎��p<��V!�9T��<��ʼ�K��i���������<=��^�O/������K��.ا�H��3��?�)|3e�_����Ê���}���_9>�4��?~Y��>�����m����}s�i��������,&� ����w�Jw�y�ѭw14�E�e��A�um��y�����2�G�Cc��ҍ<A��t����e$��̻����g���iS����Ly`)Ձ�T�Q�����������>(㻦i��O-%k�m���s��n%CI����Ɵ���� �k`/mQ�w��x�(�k�ٰ7�2*=��:�L�#�s�(k�ű��"���P��n���((?���Y���=:�{L�%�_6�ɴFY.�6��>P�Xw�𚸑}��J��C����>�����������g��6���_o.��P�}�:�ݐ멌^���K�K
K���d�>��&����\��I.K37���|���������gY޿��W{=<k���]j���������z�����NZz���4�X�����/�4���\�G����1^�V�|{��M�D����χ�>ؠ���>oS�܏K%���'���������L+F:�!z�}�߽�bx�Y}���7}����2�c��;uY��a|�^�3i곮M�l�~�j����Z�V���] �LF^pK辶zF��jğ�;�	�8�v\��:�a�{*=9����8��&k�h�v���ӧ�[':�H#ڿ��6��+[�uYP�]�8�Z6���l20��]V�h٤6�! ��[N�:��\h�O`�ML溸.������3���^���;x�~5�W��8A-�YP��V�Vʩ8��J�Pr<�q�n��3�Qd��_���Ŋ���S�{f�z�٤e�%��ׇ�7�_�?��>,uc����ai���B�������Po�6�F�3m��:ӧ]y��Mef�!�\Q���_Ѱ��_��/ҽ��{�,U�Z��x��u�04+;F��[�b5n� ��7:�u�j��H���<�����sVf�,c��=���N�h��妝��~�6=!�k ~}�mo.
�!��?�p�=|�^,U�Z�����]z7�%�����6+�����ۺ���>{��˻���������H����6�]�ލ;��!�v�縻.*���˫����g���Dq�̌����BB���Y��۫��/��F�?}��7��×��Wc�t��������^�������޸\z�2j�5{��&�5��Z�������\���dcӴH���-��%ژ[{���毭�9k���9)����֌T������]SĿo��[����n��q��Q�E���U�O�y3������m�-`y\���!ܳ_���J��ZE�߯3�F�{�e�_Ƨ��ag۲��i�3��e��1�:�6�8�L}���ԩ�7�#�`B���x4���͸H��閇��[���K6pf�F�'%��W���[v���Z���? ��qhs�@@������2�	/'oU~1xv�e�[١��KfTQc�0�5�r��]6��L���r}KYW�l��b��E��A�}����XÜk�dg�m`�?� ��߲v%��编kԽ���b�����E���ȥ�Y��=s*��83�h��A 4�?8|�ꕁ_��Z�?hu�>fK�˱ɧ�	��š��=�\ʬ�`�:��*��羕�[>�||�&GU�Yr8O=�T�YN���#x�Ab�[�����*���<ϘV���[�N�Z6�aP:th OA�iѼ�,�9�9�+��hge:���@!H#,�F��"�?��7��"^�y3�>m_,���XĤ�����[�`������&����V��2kA���!�������]�"#��[�f�	�p���r@��G�z+��t�tH�tN�J�[��;_\.����,c�%N���Ô����l/>�Q�9�s�~N�6g�byCp�k��P>m�^�i�"�6��g<�������L���9}rx@"���%�[�[�	Jt��pD:�:;l���2�5~�g�����݊���E&>	;�Ik�&>��oit��`?}-�B5�;��&p��l��Q��z	����1�zFO^3�����<�5����eB]F�&�o>�0�o6���)�׀��\F
m��ݤr?��%�[M�f�+5�q�]�X�)f������\�;k�T�0�M[1����R,$`8k'�ù��]V���3M��@2_��w,Kӵ�ݲ��9�͉K8�ksgۧ�y�ї9���J-Ǎ�ͼ��eLSU�9	�".w�(�����MR��J�b0�F+�2&�=3_�5��C�&���w�ˍF��Y䳠n��a�����k�^^�/�z-�XDf<v��|�����~�ANe�����;��.��k��8�%�%�DOv��%��"�/Y�2b&>�|�'�(��:�q����WG��]V�X���������������CwU_�_�I6q?�r����ͻ��������.���۟/~��PK
   `�tV3��Ŵ7  �;                  cirkitFile.jsonPK      =   �7    