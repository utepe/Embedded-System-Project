PK   j�tVe��D 7  V2    cirkitFile.json����6��_�Q�=��^E�b�7�]c736�s����~�[����~�{�{�#�UՙR*��������Ÿ�$�>
����xqW���ٴ�w���������;r���w����_��Ň������/w��o/���~W?|�Us��]s�l4�n�PM[�Ө��5��>��7z�/�}�����-Ao�����7�����7��+Ao,��+Ao��+AoJ6W���(�c�����7��æ��5]g�B�,��{i�m�ɷd7ႇ���[�\	:jaW�n����]}u�K6n�뻫��M��J�Sj�Ib� |=���=�]��hn�z��o<�""��`����-"R���H����)�m[D��:`⋈=M~��-B���M�u�݆�$���|�;�8�x�z|��f��nO	g.%�6|�o�.�-"Rxf��xd���SqߨB���)2���-Bo
~S�)�M[D��7El�0����&�-"R��c:���\a|#~��)�![D���l����"b߅5�S1�3�w����""�R(���X���m(�PD����l5�����%�SX舐�7%v)��҆� `*�r^�حε1w���[?�o��"ƨ�3�WBV�y��㷴��ҲED
~K�)�--[��8~��)��U����9�E[v����ibxv㹯�o��a&�y}n_��u�j։Ӯn�� ���-����FĎ�ED
~;�)��4[D���lzS��i��H�k�""dr&b�w����}���˾c���|�c��'��dt�#�D'0q���	JGX��bug�����No
��
��t����9Vw�;(a�b	�;�����t�g��]�����tz㱺�X�A�K�7VwVwP:��������t����j�۳��8y��5���|i�X��������<��f|���3$Ǿ^��V?8����/�M��`�̗vՀ�u�|�K�����;X>�L`��C,���,���a���|i�X���G`���<�_�|�K;����/X>󥽆`���W��+��À��?�|�K�,���X>��`���,����T�������|z�+)��g�k�P��Q?8|�n	f����X�Y1'8�1���G`����>�`�̗6����~�|�K����G?X>��`����W��������G`>=KD���ߌ���ʘ��Q?8x*�����|)�X��	�G`��-�?p��#0_���8|���/e(��ς�,��R��������}��r˫f�\L��U�|�|���]��}����~p���#0_ʂ�zwz{8p���ɂ',�;��r7�Zp�d�A���|)}X�	�G`����?pЄ�#0_J��8h���/%���ρ�&,��R�,���A���|)�X���G`����?p��#0_���8t���O�Rm!�A���q�9���d`���,�;;r$n!}8����/���`�̗����}�|�K����+�����|)� X���G`��3�?p��|+S Ng�͞�+>MU���4A��D������2��,�[q��N�ꭦGq�|�i�ߕŧ{W��՜w̧{��'��uh#���}|�z<�C���][~��|m�� k�3���y�k�O�\�?݅��Z����3;�r�!���H,�5;�umy��3;�tmy��cJ����﹏gyn�m4�s��X_��̵�{�m�g�RQ(;e}mUe�A���.hmZj��볊3����g_��3W�z�����K�`��ņ/}����	5����F�`F >�z�ӗ{pYŗ;pYŗ�oYŧ���?K��=�J��=>J��=�I��=>��x�z<��2�Y��:����Ы�J�����tő�@V���@YV�n
��>*�֮P������˸2vl�<=����I{L���[�G����6}oC����g?�r��f��Ee����"8�롳eW�79����̧/w�|�W^�C��:Zc�)j�+,���p>��2|Vq&�rr��:��.�Zٮ�&������/�{V�#�BD.�*���7�o��u�{k�c�LV��Gs�u;ݽM�+tmt]CPE345=y��<=���ӛjmU֪��h��U��à:[T�1���泊/?ݑ/��V����ۢV��RUрB+�>�����O���^Ϋ"��b����j�n��|�޶Ǭ.��������T�����1g��nC�M�cV�S|�隚&~�����l�FgE��wU����i}��Y�ǧ�4��<�n���ۻ�w?r: ������s>1����$H'/�!	���c�@�t
E1D A:E�"� ��THP�5����:�#�(�
�#��t��((6L� 󐣯�08f��k��6�o��o?����s�(IzE 1��7��7J�'�AL0N �K0Iz��1��8��/�$�q�Ա��q��(Iz�c1����-�����[IMSUl=��8J��$I�e2�����q��1?1��b`~�T�����q��(Iz\
�a~���q���cƄI�����̏�$���0&��t)�$�	��X%)%G�1��x��(I�
�$��a虃�0?na~%i\��X����mB�d��޷���h�L0?na~%i\��,̏[�GIJ��`L0?na~%)��M�����o�N�L_�`~�=y_�5����n��e]��e2���{�u������ok�6�F��I�?�`�q���(�����Q�RB̏�0?�����`~����,Ib��>�a�{��N���CXg{�!�z3�S���i�
�Ta%V��毀K�U��DX�f��.�W	Va�q��^�	�0�`%����4�F�$��("z�f��h@��DX�f��.�W	Va՛i>?�T�^%XI�Uo�y��R�z�`�����`� K���DhI�6�m�ѭP�%v��]$x�L�u�1T B�֚��V&��%ڴf^F�2�-�Ц��2����DhI�6�a�ѭL$&BK2�i/��ne�1Z��M{Jdt+��Вm�#�[��L��dh�����L��dh�^%���e"�$C��\��VhFLhJL&.32q����DhI�6큓ѭL\&BK2�i/��ne�2Z��M{et+��Вm�[)�[��� -b�Q�6��ѭL\&BK�i�s:F&.32q�-�Ц=�2�d�2Z��M{�et+��Вm�C-�[��L��dh�^p�
�VZ�(�2qY!��Вmڛ/�[��� -�+B�r��V&.�%ڔ+AF�2q�-�Ц�2����DhI�6宐ѭL\&BK2�)��n�L\&BK2�z��'�ne�2���W��+�Y��� -�&B�r���V&.�%ڔ�FF�B;Ʉ����eV&.��چR��|�AZ����ˬL\&BK2�)���ne�2Z��M9�dt+��Вm�E%�[��L��dhSN-�:��L��dhSn0���e"�$C�r���V&.�%ڔ�MF�2q�-�Ц�s2����DhI�6�ΓѭP���2Z�w�/R�2q���XcP��d�2'��Вm��(�[��L��dhSnI���e"�$C�rd�趔��DhI�6���ѭL\&BK2�)g��ne�2Zʣ�xFtW;k�Ϊ!�VY*zU��H'e{�i�-٥s�WJY�M�R�B6ٕR�x��bw�WJq��r+�,d�^)e!�J)�ҳ3OVJs>�^ku��Ώ�[+f����zk�`�w�ֵbRǯ�pj�Z1^:st���4�kŌV<?�e��{r���L֊ٞ1;�y��/�w�VƊ�΂\+f����k�<Y����bF+�}�V�S���ik[]LGb����b��EoJE����U�mښ���i�9ݫɒ�a9�AeI9�=yo�:4V��ke
*Q�>t�'[�*����ɒB��FYRF��O�Z)�8僳�X�^ή])�dS�%�dK�%�dC�%eᄏ�V�Oy�<1t���1��o�����3��x��bN�+V�Ψf(��.B�**]�TG��t�i�%��-���MaU�Ƿ��+Tp���.�7�26/�Y���d!�m0UTj�!Ji�jU�WC������Y���n�\�z�P�ȚF�EpJ�Cgˮ���QGYR0,'[H_���W�����B���;E�u��PuN�Q���o�%�F'��!4���	�r���ڠjr�czj��κ�zɒr���sC��QVU���k�UoT�����t_c���,��u�Q�M�.tmtvCPE345=y�O�dI9��TCh��VEU�/ �J�uTg��4�#�g�Q���,�|�U�RD}���
Ɨ����huNeI9�2U=�WE0!AUC�*�-�.Խm3l7G�i������T������I���6��}�e�n���,��&z�NE�YF�з�cRl��*U���,)�,?�b6�������x��G��K|7���]}�˷��1���w
!	�c!	�c{!	�c\!	�c�!	�c�!	�c�	!	�c!	�cL!	����"q^�a~�`�%Io�0L0�M0獒��&��&�GI�ۉ6̇̉�$�� �	��̏�$���$�	���u�a~���8J����b�`~���8J���c�`~���8J���[c�`~���8J��Ψc�q�/`~%)墄1�FRpC)0?^��8JR�c�����Q�R�:̏0?���r���`~���8JR��c��q��(I)��	7&���q��(I)7�	��-̏�$�\00&��0?���r���~`~���8JR�uc��q��(I)��	7���ބ�q��(Ii<�	��̏�$�=�0&�/a~%)��1��x	��K���ם�GK�n�H%Va՛�^p�T�^%XI�Uof���R�z�`%V����BK�U��DXc�%��YZ.�$XI�5��D�:K�р+���>��^g� �`%V����BK�U��DX�f��-�W	Va՛Y.�T�^%XI�5�	�	d".Z��Mk�et+u	�]2q�^$y�ВmZk.�[��K��dhӚy��D`"�$C�����V&
�%ڴ�AF�2��-�Ц�2����DhI�6�)�ѭLD&BK2�io��ne�2Z��M{|d&d�2Z��M{�dt+��Вm�s%�[�1�)1�����eF&.�%ڴNF�2q�-�Ц�|2����DhI�6�I�ѭL\&BK2�io��ne�2Z��M{Det+��Вm��*�[��L��dhӞ]��I2q�-�Ц��2����DhI�6�ѭL\&BK2�i/��n�V+
-W���
������DhI�6�͗ѭL\&BK2�)ǀ�ne�2Z��M�dt+��Вm�� �[��L��dhS�
���e"�$C�rp�����e"�$C�r���V&.�%ڔEF�2q�-�Ц�.2����DhI�6娑ѭ�N2��d2q���ˬL\&BK2�)g��ne�2Z��M��dt+��Вm��$�[��L��dhS.*���e"�$C�rj�����e"�$C�r���V&.�%ڔ�LF�2q�-�Ц\m2����DhI�6圓ѭL\&BK2�)w��n��|����˜L\�d�2Z��M�et+��Вm��(�[��L��dhSnI���e"�$C�rd�趔��DhI�6���ѭL\&BK2�)g��ne�2Zʣ�xTtW;k�Ϊ!�VY*zU��H�i{�i�-٥s�WJY�M�R�B6ٕR�x����y{���\�+�,d�^)e!�J)�WJY�����@Ƌ�ޥC_׊����Ѫk�`,x� ӵb06�tL�Z1+6+^:?s��/�R�VƊ�΂\+c�K'.����s׶�+^:=𣘶q�3M�(��������B[S�6-5�{5YR0,'?�,)'�'��P�ƪ>x�lCA�"jۇn�d��T�i�dI9��,)'��%���n&K�I/�%夓ɒr��dI9�b����0yV2^�����������^���lu��j�"��"���ҥHu��MW��2YRN�SYV�n
��>���]���Uw!ĸٕ�y9͒%�$io���R�QJ�U�R�ڦ�m�?͒%�t��Zo�Ы���F�4�.�S�:[vu|��:ʒ�a9�)�qE�U;4>�Ъi�NQc]a)T���-G�i�#�F'}��u��t9��vmP5��1=�ASg�i�dI9]�޹!��(�*J���7�o��u�n���1K�I��	ٺ����&g�6:�!�������קY���di�!�UY����\��:��Eeӑ�3�(K�IG��*[)�>Ji�Z�KUE�M��:�����d���׫"�������j�n��|�޶��#���v�zW��NY��Фv��N�����.�vs��d��4�;t*z�2z����b��U1�*�uK��]��.��/q{}{����v���ˋ����͇�::���������.�}�5'�du���d<����X���N+��%���z�fET�G;���d���Hfg�푰���٫�֌���y0����Ew�9*�R�t+�Y�[�=;=��r�9����7����^�.��?�ۗ��w�}�(A�����b�-���{<�S�|��=�2���\���<���u�8�����}<��+��Z�����1���yL�gy.���e��]f�Y��qN��}w�&�WB�(��B��r�2Vg�Y)��f�z��,�˳���ܹ\�tSK54���	����ʅ�ɜye)bz���(�̕/��_�z[&�י�R��Y&�]~�$av����%^]l�9fd�=���3>�
���I�3p<��b�!�V��j�4�t�&�u!;)�J�w]�:8Og�������>�3�x<���C�6�=¶�2ᜇ��x���x
'���NűU�������ۿ�ݦ��-��:�Ǜ�����+� ܅O ��' w ���O ^��@�Q�>�%R#�SO��U��ז z�%f�Z|} D�qW�%x�Ep|"�Z8>`IܲW\Op�¬n�矴�b�!���W�XmdϏ���]���n�[������WX��tU�a>S������x;v�{]O�����`��<��R/�ZZ�{6���X�� ,�P Vf( �1��]�����P_*w�8���vP#lT�p��H���e� ��_�· ,r蜷�1����g��O`<`8���̉X�U� ���g����v̗�ݵ�� o^xe��)�O`+�À��p�ҏO`�h+����hm��6>z7`%��ƃ=K�q�s�ʃ�'��_��/��l��Pq�� &� �q � �ʑ���n��h�Nk�&��^߭��Į.|s�
��K��_a��@�rގ1��P��;�;��&��3����)4p�ss#Ɓ0�8B��VG���G �	���O�F,E{�p	�-��*�enH}�� j��9�����C+M�J;�0�vZ��"��X2TȺ�lE�X���������~�/޽�~;�'ln7�W�Ż9�t:=a�Cf�؞¤`���I5L
�=�tä`���)pL
�=�"Ǥ`���)tL
�=�b���QŃ�|����=����>� �iz^a��h���B�Z�����3� ޗ �/CoO1�r <0\0_�ޞ��� xab;M���s�� �KlOI z{r8��p��^�2���r.��E�"qp���	sR� �-_��ξ�j�����"�X �˗����O��	`ڊ�bUs,Vڊ�b\3_Fh��/#r \3_F� �f��ȁi tu�����i��1w���!� 8_������eD@ϗ/#r �+_�8�=39֢ڊ�b�-_Ƹyc֥b��Y���N�f�Yİ��we�)s ��\3_Ƹ��?� �l��/#r \3_F� �f��q��/_Ƙ(ef�����"�X\3��8�kv\3�Au ���Y�Fch+��u`Ȃ�����D�eD���ˈ O͗9 ��/CoJ���ˈ�^3_F� �Q�e��s��k��,��̑1Wi����}c�����̺�).K��̷��?����|zS��W����#0_�����`�a���&`�9���|�}��J���|��֟��G`>����������O����/����e68�����,���g�nKHh´x�CxP�J�a�4�
T F�3�I���j N���*E�*`BB��h��0!�	�bm��1��Єz/�F��L8O&�et�B��LHh´��Ct�&$4aڜ��!:��0m�@c��0!�	�,�%T F��L�gI��1:�O�����S:N�0mB���		M��9�u��S���&L{��:D�)`BB�YzK�@�g���0�
0���c�Q):l�S��x��Q�AG1`BB�=���$�(LHh´�Ct&$4a����!:��0�[E��2�4��(�@G1`BB�Y�?�@�g��%����i�3Z��LHh´O�CtP&$4a�c��!:��0�G���		M����uh�a��Єz��N��a�p~\�lgk��h�W):��N4�<���A�U�j���&L�+�:�oy��yA5�LO��2zjfN8�e����U�j���&LN�:D5`BB��,h��0!�	Sf��A��Є)+X�Ԁ		M�2��u�j���&L��:DG1`BB�\Ih��0!�	Sb'��a��Є)Z����'�b�9N)��*E�-`B:@8����t��Q��Є)sZ��(LHhu�Ct&$4a��a��b���&L���:DG1`BB�L}h��0!�"\y0�,k��#���gYW����]Y�@�o�9����q���+��r��>��xr�է ?�q����OhZ|�������(��f)��
���_+�k�����
�%�]+���rg7s��O��V��l���\�=ӧs�v~��Z\�5�:ขgwi��=��xf3�q�q����
8ұh78Ӕ�B�)�k�*�*�5u!�����d��>��G�U��7���X���m(�PD}���l5���p2�!��
Mw��g,��,qE���w�S��qe�;u��JqGZԬ�GԬ�G�Ӭ��kM�i/��<yl�c=�v^��y��ֽ���8J�q�8�b�>��u�Q�PD�_�^UT���+�y��G<wYV�n
��>���]���Uw!� ە�!:����G�O��`����C,�z�8������{��=?����˵ޚ�W��ߚF�EpJ�Cgˮ�/sT�Y��?�r��5�(�j����/�jھS�XWX
UG�V�#�Y��GZ�!4��h��je�6��\���ڠ�����g�?V޹!D겪by_��z����]���;��d�?��h���b�������h�h����'����g�?���B[��*�:�op���0���iLG�?����G��ȗ]e+E���mQ�`|��hI��u[�V�#�����ϫ"��:�AUC�*�-�.Խm��_N�c��ۡ�]�Z?8e]C���;݆������S���55M��;}X�߾���b#�U��^UN���*�}�O��]u���Mx��ǋ� ������:������L}�L�@���^��W{�����x��c�1�Ƙtv��L*1�n�(ٸ�Ҥ&�0��I%L*Q�1��&�VF�3Ǐsz#������l||\,��;�+�Ӝ��i?�5�Ԗ���wNk������
���9t�@���+���_:ç��q;�#x�~�7�C��7�b��o���-XSR��Q��D��E�ދ�u�)'�g��^r��;�����5�2z���h��c�.���!���58��垿��g�kiL!w|{�:��:�Q{����6�������ۅ�&*sĘ�<m1"���{f�,0g"�z��o����9t��g�;��3��Sw��j����o�
N5�r��W��x�;��d�:�9�g���a愁KȚ��9�����SY8eu܎�a�S��М�\B�A�L��:�vu-��tV����s�����j)�7����I�����ŀs�~�7F�1	�|y��������:���s����?�oR<<�d�.�����R1���.��%z�D�K�钙_rO���R�t��_
O���=��^0��k~^������+�+��ULs������ߎ�g�_�x�g]�\��l	47�3W�y������w7����h^{�Y/�h����f�#��n7�W��Pc�Q����c��w�������?��u?<�c����gt���C����/�n?�wW�8��݇��������n���M�]�=]���k}��~�MRi�j���*�_ğ�����F������������j��������xu�w��Ī���y����;�{��]�xus �(�K^=\�F=|�|U��vG��eԹ��L����.L�5��By��V��ֱ⪦����q������i�e���./n�bu�[����O��]{�?U�ת�����U$��������]��r�4�R�b�-��%J��z�����T�,���.,��J��sZ���r�b�
�^�;W|UN������n��]*a�J̔�t�����|aV�f��|aV�f��|aVO浐.���K߲���p{��w�?������_��G��~������U7���Аv�j�`�-�����+}Sն����>\�F���]��l���R����m�U]�ta��D����lz�N9�����R�!�l��;O���L[�Ͻr�K���|x|�)l�ֹ�T_�YށZA:����To_��w7꓈?D���U���^]w;�۔>�z��QrtDu�uј����ֽ�T��������͎�0�.��U�D�d�jPU5tj��wu�w@�o�o��]mzO�%E��Jj�^U��U�)��:O��/�P�t}*��o�[�u埥����lnF��ݻW��lO�������7}y{�𛮻����tI�ָ���?`Xoc�]�o+��R+[U�걶���{jL���k(L54Q��o�lf˶�U�Fôֻ�����r���j�!>�z\�c��hr�Хn���)�&V^WW��kJUuu�8:S4�@]h����n}��۫��}������7?����?�ӛ��7?�>�m��Iw�����/�<ܾ�{�ys[�w����?m�3
���=,���怘��C_?����¶�_��}�0��H�ӥ���z�ߧ8�ˣM�M�>���q����cwu�o����q���VG#������?*r��@����|�x�������'_V&6��p�^߈�"~5]�K�y�Qt�U�=mtw�_�E��ӾQ�Z�iߨ���f�;2լ���l� c��e�|�xn�Қ������Ak����}c�WY�,���8�73��0��Ķ�������n��T����Z��C��Ի���PE[+��OudvM.��/�bP��+�2��ұ����t��lƸp��VQetǣ�}�*�~��g��x�K�s5���M4��;�oX<_0;7��^,��۹iү��¤'�r���_.���F/�N㆗������}���/�4���?|���|��gw�u_O{Ke�/6�>F1�2/����T��ף�n��]S��ȶ�]�a�}E][�q<k��Z�飋}c��ҍq�I��W�\F�ϼS���?���/m*SC1�UQ�YJ�g)U�(kj�ilPu����*6�.|�4m����d- Ͳ�ql���ѭd(�}�<��篾�2v�y�׶�(����M���ٰ5�2*=oM���Z�]�(k�Ŷ�+W1������4��;
�e����Y���=&��6�ɰFY�ml%}����́�č��?UZ���co����>[����o~�2z����&|����v��;���\Oe��U>���~������G�҄0sCY�3zxa�
�e17�w�0�+���^��8�����_m��S���c���j߹�ҍ�/����臘Ǳ�I��%��?�7I+��e��|t�Y�����o���)M~���x>����?������~�*yk�?鷴������I���U�c��8`��/䏏�5�ݛ/�7��7��Q��/�n�^�Z�z���?�K���ho�>�4�Yׅ�6Z�s�K���Z�V���&��/ ���4� ۟5ƿc� 2lc��s�c�cH<�����)r��St�{[E�>��&��O��^����g�X���5臺TT{�}�"6�3�lP/k[WV��؏
Mq�+G~z�3����86�Q�;��@���d̊��6N|\�13�9l�7��elm�.����^�
�@k�@L�fb|k�[�����%���6�f��c��p�
�ʯV��bŊF��qj�����Y;�s[c$4}��}����g*�vKݘ��l�T:9��7L=4�/�/TMC5E1��
}쩺�O��?����9��gf;�a`���_�{��vY��6U����cwC�2/���V��46�幋~��_��k[v��qovÜ��#�X�s���X'� ��r�r�
���g��~HW���Oöw�b����_uߦK]�5����o���|��ij)}�����a�Q�m�~�w�����x��߮���=V�ho?�{׷w㊽���s\%|�����Ӻ���lW7�tDqS������B�Fy�"G����������Q���߿�H�6��L��H���N�;���hy_�~@��C�U�>x��[1�}�^��4�o���?E��%��4�Χmci�6�n۷��mK6F�ڣ6vNz�#v�6��)��������g}���b]iU�ˎQ��F5��
�~�f&��_�[�k`y\��
�]��_w|�^H�}[Eo_��n�������/�3�ڰ�mY������e��YmX��m�`k2�I��Wx�N�����6���	��m�I���;ܜL��mN^��3��V0�9)�МL��qc���� �5m.�H�\��Y�B9���]�?��٣�����KfvMQc�0�%߲�=lR����������L٢ͥ �#h.ڷ��̥��kg�5^��3�ӊV0�T�
^��wY�Љ��ܖ�ר{ߣ���A!h.��
.��װge�^g�w�`�?�
^��wY���sn����ڧ�'@s96��:����8�?�g�K��?�̎-D{{�s���-�>^�#U�Qrx�z��l�7�2��]F��	b�]��������Ήf	�3��fjr��ӻ�0h:� O��Ӣ�γ��1��i_Q�vVEW���-0�#,:�8+�S����pV�՛y��h�b�:+��Tݒ{޿��2��M�-�ɾmi��*�&��o[1���+��l�����k+��p w��:/\��p�r{�G��uW�:-��h�鐤�h�0�k��;ѿ�<pWnugDkV����^�*���̈b�՝��s2�9�)/μ��"�O�x��M}��s����'���m������(�vq��/p�D���x���!�偻�-�9G�a���,�^��~�<o��-�y_���'a>���$���C�k[S�L�Oo�5�P�ӊ*�	DV��'X�={�Dɘ0=��'�{�w��<�6���'1B]FX�M8�|�a@_mLY{S��-�9�Z��s/� >n��ך��r'Vj�sD���>C|� ��5 ���Y����a@/ڲ���N�?N�B:g-�b���*��]󑦃�@2o��w6��k��d+����>�8�ssgmۦ����ǐ��*}��8Y̛y[��4U�0�%�r��'ؽ���h��eS����0ZH�1Y�y[���n:t {�;��<j��ȟڋ|��xc����xz[eO�gݖk,"#�vĳ��F<�Nx�J���\�=y�)���������x�,�~�������������~���������.~��PK
   j�tVe��D 7  V2                  cirkitFile.jsonPK      =   -7    