PK   -�mVRe��1  ��    cirkitFile.json��r$���_e�{qA�"@�0�Y��8�RX>�Eh���0E��%�Bt/s�t@5����F1�)�k�nX$����D"�, ���n��W������������:{G���C}�}_��U��}����]o�rS�p�������c������Xf��t[wF5me�-�F5uݨ�p>P��z�7���7ߞ?_�%�����`3p%�a3p%�e3p%�c3p%�M�f�J��f�JЛ�����7����}�Q�ED
����J�;K��H�w�l���0�""�e�ED
��d��|��)���-"R�]'[D[�}'[D���N��Hh�}g���l���;�""�w�ED
��d��|��)���-"R�}'[D�	���-"R�}'[D���N��H�����}'[D���N��H���l���;�""�w�ED
��d�����l���;�""Er|����}����6�C��൲Lg����VCQ�:�y�����uS_\f���ח���ݏ���S|nG� �i-��nu~*���]�y�U�L�꾈�z�i�-�2ߞ��X~��)ʅ:��c�hVBV��e[�z[�e���^�����Ζ]\o����*-��d�����-"R�J��q���-"R�E��E��,��v�>�^=F����wʎ�)S�y�����.ݱ�t����Ow�I_�z}�}��ǯ�:��Fm�CZ��H���""��f���~�-BoJ~?�)�!-[D����X��u���f���0�U��c�Ы�	����2�	L���xz���No
��
��t����՝��JGX��cug�����.����sX�A�KG6XݕX�A�K�7�;�����tzSauWau�#,����VwP:�ҥ�����l���B�̗������.��8� p�A��G`���?p���#0_�D �8����/m �m`�̗6n���8�|�K[N��GX>��2`��#,���6�������|i��38����/m��`�� ߡi���x�9�T��FГ#3�g���s��WK����G=X>��`���,����E���Q���|i�%X��G`��Y�?pԃ�#0_��
�8����/m���`�̗������,��Ҧh���Q���|i;7X���G`���?��.��.p�a���X>���`���,��R��������|)�X���G`��*�?p���#0_Jr�8����/����ς�,��Rb��������J��.ʝu�&4a����>I{V������G>X>��1`��w�����#�|,8�����g{^�&W�,8h���/���4a�̗�����|�K���MX>�DMX�9pЄ�#0_J1�8h���/���`�̗�\��]�|�KY����.X>��Y�*�<��f|��r1f���@�_8|����gG���������>X>�<l`��C,��R9�������|)�V%8����/e���`�̗���}�|t�oe��i�ɵY�yŧiW�&�]�Đ�Zv�WXF7��x+n�܉wC�U��x�i�ܕŧ�nW���]Y|�_vm#�6Rf+�
��<����\[~z����L�[��<��ƣ"Y,�������xnŴ�ف�k�3�v���x��U}��������x�z<��:VӝQ���r�k7��)��S��VU�Thk��EK͑�iVq�ӗ~V��v���7��.�c�ׁ/5��c��O_j��gr	����r�F�`F�z�/���/����/���/��s�@�s0�s�s��s�a>ޱ�>~��q@VﺮP�`�0zUQ钰��92�*~d0�ڕ�U�3.eb�_OQlך�itul(�S|��eYٺ1V�>V���Q������*]�UG��U|�餽E�>���^5�*嫡m�ކ`�#O�*~D�y��x&8�
�@!.ʑWW)���p�x���Ujt��w�댥Pu�XDV�e��*�<0�*�<0B���>D�C�b��&����S[uT��U��rn���X��7���P}kz�E'�t�<AV���Vl�.F2�M�A�C3CP�������G��U|��M5��*ke�:�|p���0�Κ�h��lL�Yŗ��ȗ]e+E��⭩U(|��h@!�o_�|V���?��7wכ�������O�6���E��v�ӯ_�4V0�$H'_�!	���`�@�t�21D A:�"� �PH�N1-�$H�0C�S�!	�c0r�8��s�0�M0Ǎ���o &��&��FI��W�́�$�qb���s�(Iz��1��x��(Iz��1��߸8̏0?����i~̏0?����� &�/`~%I�@L0?^��8J��8��q�70?����xp_Rp�R`~���8JR��c��q��(I)� �	��̏�$��x0&��0?���2���`~܎���/ L0?nG�;��	�M|��ee:�0�`~���8J�8�<J"ߓ�����Q�RB!̏[�GIJ�o`S?0?�F���-�8�w��w�c2����oYWE�2�`~�=xߺ�=�	7�9z߶��00��7O+`���̏�$��0&�w0?���v��&�a~����Q��nsӂ$�f���x�{9���&l�l4�Uo��0�5M���J"�$ª7�p�@�J����Ls����*�J"�1���4#F�$��A"z����h@��DX�ED��tH����L����*�J"�z3M8�
ԫ+����4\*P��$�����DhI�6�m�ѭP�%v��]$x�L�%BK2�i���ne�/Z��Mk�et+��ВmZ�/�[�(L��dh���Db"�$C��b��V&�%ڴ�DF�2�-�Ц�12����DhI�6��X���DhI�V�eeA�V&.�����3N�̠t+4#6�EL�Ц�c2����DhI�6큓ѭL\&BK2�i/��ne�2Z��M{et+��Вm�[)�[��L��dh�Q���e"�$C�����V&.�%ڴgWfa�L\&BK2�iﱌne�2Z��M{�et+��Вm�.�[�ՊB�e�2#���L��dh��|���e"�$C�r��V&.�%ڔ+AF�2q�-�Ц�2����DhI�6宐ѭL\&BK2�)��n�L\&BK2�z�8'�ne�2���V��2+�Y��� -b�L�6�v�ѭL\&BK2�)G��n�v�	m%��ˬL\6=����� -����eV&.�%ڔ�HF�2q�-�ЦN2����DhI�6墒ѭL\&BK2�)���n�L\&BK2�)7��ne�2Z��M9�dt+��Вm��&�[��L��dhS�9���e"�$C�r���V(�ǜ�F�V�֋ԭL\&B;?��:�����e"�$C�r2��V&.�%ڔ[RF�2q�-�Ц�"�-e�2Z��M�>et+��Вm�Y*�[��L���h?����]g�B�,�^�}�k�m�ɷd��a^)e!7�J)�dWJY��R�=<p^)�˭����z���|�+�,d�^)e!��Z�/�z�}]+c�KG���pj�Z1^:st��oO���ײ��=X��8��b@>c�K�T���⥳ ׊�x~(�Z1V<=Gc��ъ�G_������U��u1�x���Ob���hJE����U�mښ��u�RszT�%�r�AeI9ٞ�/�:4V��ke
*��m������*��<ɒB��FYRF��O�Z)Ŝ��YR,D/�#ϒr��̒r��̒r��̒rr��gu����C��o�����cNy�<1�Ϗ�Y+�d�bu��
�&�nzUQ�R�:��EgN{�,)����jW�V�θءD!FҊ�`��tM���� G�I���l��L5kkgTp���.�û2vu�Y���d!�m(�X��(���qT)_m��6۟fɒr��\�m1���2��-U�����Ζ]_Ϝ��앲�'}�ig�W�����U�����:c)T���͒rR�YRN�?�����^��ˡV��U�K{詍M���^��dx�ߣ��(��ת��P}kz�E��t�1K�I�؄l��1]o��]�4f�4C�Qӓ��4K���,M5��*ke�:���*U�aP�5U��>�����dq�ˮ��"꣔��*�TU�����s�(K�.�ϣ�������������I�����UwS_��?I$hk"� =�H�}�$H���$H���$H�q�$H�1�$H���$H���$Ho�H���ym�ۆ�m�9n�$��1L0�M0獒���<�	�	��Q��vB	���s�(Iz;Յa�����Q��vÄ��0?^��8J���5b�`~���q�$���0��x��(Iz;?�a�����Q��v�������q���sƄ���������Q�Rn<̏�GIJ��`L0?n`~%)���1�����q���k
�����Q�Rn#�8�8̏[�GIJ9h`L0?na~%)�<�1�����q���c6�����Q�RN̏;�GIJ9`L��M��&̏;�GIJ{�aL0?�`~%)�-�1��x	��(Ii/+�	��K�_��~_�l�3Z�v�(@*�������<���*�J"�z3�
ԫ+����,Z*P��$��.���OA4 �J"�q$��Y�)�$XI�5�QD�:K;р+����,�Z*P��$ª7�|Sh�@�J�����rM���*�J"�iM�L` q�ВmZ�,�[��K(쒉�H&�"��K��dh�Zs��D_"�$C�����V&�%ڴ�_F�2Q�-�Ц=2����DhI�6�ŐѭL4&BK2�iO��ne"2Z��M{cdt+��Вm��#3� ��Вmګ$�[��L��dhӞ+�
͈	M���e�L\V��e"�$C�����V&.�%ڴ�OF�2q�-�Ц=�2����DhI�6�ѭL\&BK2�i���ne�2Z��M{]et+��Вmڳ+�0I&.�%ڴ�XF�2q�-�Ц=�2����DhI�6��ѭ�jE��2q���ˌL\&BK2�io��ne�2Z��M9dt+��Вmʕ �[��L��dhS����e"�$C�rW��V&.�%ڔ�CD�V&.�%ڔKDF�2q�-�Ц�(2����DhI�6�v�ѭL\&BK2�)G��n�v�	m%��ˬL\fe�2Z��M9�dt+��Вm�}$�[��L��dhS'���e"�$C�rQ��V&.�%ڔSKD�N&.�%ڔLF�2q�-�Цg2����DhI�6�j�ѭL\&BK2�)県ne�2Z��M��dt+��C(͇L\�d�2'��Вm�e(�[��L��dhSNF���e"�$C�rK��V&.�%ڔ#SD��L\&BK2�)ק�ne�2Z��M9Ket+���R����٢�Bh�%ӫ�/�|m��4����9�+�,�])e!��J)y�WJYȼ�R�B��R�[�����z����+�,�|^ku ��X�ҡ�k�`�w�hյb0�t��Z1^:&t��+^:?s��/�R�VƊ�΂\+c�K'.����s���+^:=𓘶q�+�RQ(;e}mUe�A���.h]�Ԝ�dI���lPYRN�'�U}�Zن�
&jۇn�d�����zɒrR/YRN�%K
F/'�L���^&K�I'�%夏ɒr��dI9�a�d��==�����ӣ�<1'-���]��Lt�&���ҥHu��Μ�2YRN{__ծ��
�q�C�B����v��FW=A���,eYٺ1V�>j��Ψ��A�]1�we��N�dI9�B��PT���QJ�U�R�ڦ�m�?͒%�t���b�UCe|#[4�6�)]�-�:�^��dI���n֦-�1^�C�^�VM�w�댥Pu2��)�=U����SCh�ױ9�r�Ul:A��R�zjc��;��,)���!��(�*J���/Tߚ�uѻ4]Fk̒r�%6![wqL���xC=��2��t���>͒%�$KS���Z���- �J�uTgMU4EG�Ϩ�,)'Y���l���(�5�
�/U�/D���:ʒ����y��X�ח�7��wT��}q��n>^���7W�뛮�9{��7���5,�����7�a=��g�g���%�ٚ9p�x� �I�#����G�~/��fd/V[3�g��΃)pj!��\t���?K	�-+f}Lw&qP���Y�t�����+��$�:i���B?���}ɫxGܷ�$F� ��/�r�~���1��-���xv�s���<����>�q؏�/�xV�W,�g�8)���1���yL�gy.���e���.s�,4�xN��}w�f�B�(��B��r�2�`�Y)�/+��ɳ<.�B�,���Y�X��oX�����}Kȿf΅-TL�KӃJ8(�D9f�|q05�z�o'Zn����w���;4��M|�x�?�_p�	���� p� ��( sV�O ��za�����5U5���{�p�W]��; ��S}�Z|y D�qg!���d$�='�'LM.{��Ϙ ;���g-�Q"�6�B�j#�;���ŵ �? �������L]��d:�U�B��0��T�;�^��=�ˌ6�D���"{�������f�+��b/���kb ��1 
�
 `��:��e��>>��r�`(�kx 5�F@�wA�+h#�_ ������A�yk�0�s�hxƘ!y� �3�H�O^\�9˾�R-�Z8���>/�lӲ�����>���^(kJ�,)�+˞���,@�esס��Y��'B�J�D_ �k�<NBr�Ty�1�Jm�}h��������/��7�w�]�����a�j`sw���������y)yņ7��M
¤`��c&[���0)�"��l�I���duL
�=&�cR�E�1Y��-B����lzL�Ǥ`���d\����	�p�|z�����p�|z�1���p�|z�����p�|z�#������e�m�r.b<���i�|z�h������e�m�w.�� ʗ���� Z �)_�ަ�熒 j ��/#r �)_F�@�� j ��/#r �)_F� �S����|��O�2"���e��S��q"���6�B���bbܫ5s,��ڊ�b�q7� ��8_��q�uVk������b�����|����2��|1_Ƹ�`f�������:�����\�;��YK^i+��5w͚���"�Xn���UL�D��I F�|��w �S;����HG�8 ��xj��tD5���K�W���
ə[`�u���9��#~��K?K���כٱ�̺��gΒG`>��U��ovf9�}�|��֟��G`���g�����/�M��s`�a���`��`�a�̧7�?����|zS��W����#0����XX>󥕗��l���b		M�V��u�B�a:!t B�HLHh´Z�Ct4&$4aZi��!:"�0��F���		M�Vx�u��L���&L���:DG'`BB���h�#0!�	Ӯ ��Q
��ЄiG�C5:N�P϶Cbt��S愓�-f���&x�J�(3�Ӈ`�G�Rt&$4a�߃�!:��0�MB�ŀ		M��U�u��b���&L{��:DG1`BB��lh��0!�	�^<��Q��Єi!z�:��0�D�ŀ		M��o�u�[���&L{O�:����/�B�)�t�&$4a���!:N�0�WF���		M��Z�u��S���&L���:D�)`BB�=�h��0!�	��|�-:N�P�%�����	�9�g�}<S�ŢÖ9�DN>�J�Q�EG1`BB���!||:���(fz�
���Q̜p23�:1 �A�Ԁ		M����u�j���&L	W�:D5`BB�d1h��0!�	S��:��0%�A�Ԁ		M�2
�u��b���&L��:D�-`BB�\Mh��0!�	���4�@�g�ǒV��cT�[���U�[愓:2L����b���&L���:DG1`BB�Djh��0!�	S8�Kt&$4aJ`��!:��0%�C�ŀ	���c�g�מV�,?K|���,[��c���\)�@�ׅC����Ҩ�,?K���,m���t�k��m�\���_�V �B�'ƭ0��V �燫��5��8�I;�����r��(�N�z�����Zk8r�p���<��Tsyđ77j���gC�pĊ���hJE����U�mښ��[j��F��s��e�?҆�/�:4V��ke
*��O������*7��g�;p�A�w���g�]r��#��ƕ%��Hn��g�;҅f�?҃f�?ҁf�?2��3��������m�����ͭ{�7��;p����;pp�B}X��B5��߄^UT����Eg�y���<��jW�V�θ��Ģ!�mEu�]k����ў#����ee��Xe��J[;���Uw!��ܕ�#<����G�O��PT���|�U�R�ڦ�m�?�������Zo��W�����MpJ�Cgˮ�/c�\�`�Y�歛��,q��37m���e�jھS�Xg,���pL�Y�(;���aJV�#Ô!4���Nu9�*���jr��=���t�{���G�sC��eU��>�D]���[ӻ.���;�ز�y~l'���ஷ�y�.�3e�����{}��Y�<����Ve�LUGs�Ru�YSMё��?����;�eW�J��|kj
_�*ZR�������U~�����>���6wכ(����Og9��ٻo�R��z�Գ��+5��v��H�4�MC�q`9ǯ{cO7N9�Njt-��T�R�"�(F٩D�J�D�J�D�J�D�J�T"F@���ʈ���`N׍z��������ҋet�{r���9��>R���WY�s��<XA9�m����h�@��+����
�4ѝ���o[�U��&^�b&��h���lΚ��̱&�&��/j�^�Ycr�R�7K�j�	�Ԅc}��1����h���;�.���!���s�w�ا�_�����Rh���v�:��:��� ��~�e��`��q�va�{���y�Ҍ���X�=s̙�3G�̵��l���:ͤ�tTpFNL�MI�FN� N5�r��W���x;��d��9�[P`�:�4��n)���ǣ�v ��������e���)x�x�4-���MLN.هKv~�<\2�K�ᒞ_��K4�T<\*���%7�T=\���å0�D��4G�'���᚟{ħ9?=��ʢG�\����4qz���C����r��Z/����������OÛ͟n��M��m����O�Rl.��n�_��O�����]������n�?�7w���컏W�?�)EE���\\�����.���������O��*)�L�u���O�������(���P_����m��ۋ���M���7}w��.�G������n��o��c ����t�W� ��}����u��7�W�[ow�y^F������X�0]�6�;����U���V5&��;o������]}�n�d}�<?�����Uoa��?�?�7�e�P�ߨJ����W�(b����e�p�.�0K%h��^(Q�����.إ�R	Z(��B����8����-w~1�Wh��޹�r�<-\pK%�R�b��L��j���f��xaV�f��xaV�f��pa^��蟺Ԗ��·�ˮ�9�����ߟ�{v�����������E7���Аv�j�`�-����	�;sSն���/�������.�P�kuoR��
e���q�@J�����vuaƲ��;��{��Ju9e���<}�-�h���+�?���������E�:7t��M��?P���BE���5�������$��Q'�}է7����e�#�ئ����u�G���]�Ec*lW�������뛛�/?�W;R�@�,�Z5MtH�T����S�������)�_^���4��=u��>*��{UծRG�2Š�����c}���\r��o�֕���/���%�w�^�ãY<x�7��_������ݯ��}��9�Gm����z�W|�X)E��)c\Q�*z�X�V׍�=5E���k0E54Q��oKe�*�m�V6��ޙ>2�:��E�U3�Iu��X�>��5��͢q�+ʪ����U,�RU]GW���m{ܸ�����v}ѽ����?�������޼��{�������7��7�����������7ױw{�����?������r��/����?��]�]��+lK�uٷwO���>?�:�ߥA�WG{n��}�@�zq���}wq����v۷�[z���p�D_����+�+}������W�QQG
�*MU��BWѝ�ָ�v�;8���f�E��WE?[�q��FVm�����f@sG�����i��wF�t!�!������}'z��\-⿇L4����ߊ[U�
l�W�7����{�۫�>��o��e��{������<Tq�e�Օ��X(��l͠�W�T�KǮ�n���r1N���X�dy��E�M�
idCe�����_����?�����;�oh/;7�Ǜ��?^p;7MFr�>^����.��h��M��t��t�4Rx�P�=������a�W��Ϳ���_)#�W�t>�����:xwlI��b��s
�m�c{Գ�m(U�yC����A(��b[�A�0辢�-���^C�Z��m2�G�kG#t��!+p�r���V_p�����dO1��04�7���8�7с�U�^?��i�1x?�s���X�q3�`f�4��\�e��W�y�����_��6�",�ʣ�=S����55�hlP��U�U���X�m����d���1�",�JQ������/�2TX�
�$��P��7�������z�UT�Q�GY�.�ͼr�P(��A�mѨ��(h?�q�2�#9�r���q�_�_����_>g�X銸q|���K���Ӫx�/�~6����o>��/`+����fC�"5���ߪ}�z*c�S���,�3c_�{et�s��hB����e�&S�D�v1~�<t�n���U%]���?�o/�o�S���}����ݹ�v#�S����;���ڤ�ƒ�뫿�հ�<�ԞB(��q�(��������D�����O<���dl�_S-|Lp;�h�-�?鷴�����s��g����4Cu�gM���5�͛/�7��W��Q��O�nў��2���v_��lho.�i�n�$]�Fim:�\k���j]=5�E�9�=��#��m��1��#Ulc�Z�m�#Ѓ1���i�� �X��.�Ƙ�� �ǯj#���k��/�������V,�$����q��+���)�ܵ�6	��vP�X�~�KEu�T��@��]��&���L����'�k��wH*�}��ā�7���嬝��O_��}ٸ���Ͷ�w��|�~"p=]�ְ���뺦>��zn�^��x������8������Z0��g�e���a����wS�|>w��n;e�i����c�\LW(^I�"��ߝ)҅~����݇tc���E�!��C��ސ��L���ì�{H����C�}��Z�������?_���G���2J+7.�oƥ�A|�q�D����WWD���r���; ��Er}S�55�����닫�����޿��~9|�.|=�n�_�}��w\<��7�ro?e����mqHu�6�7��}~�-��}������]�=��tK�붱���6�l���o[�1�c�6����G�l�n�Sv�	O��7*�}�)e���=�u�U�Q�Q��f0��
ӻ^_���Y�^�[�+X��[n��3�*��cJ��m��V2�#���5�5�Lk�g`��;�О+ɾ����>3��F{ͻ-��e|�:�6`�s��H���;"z���lw��pO4�+�'z�
�LV"Z�`�R"*��w��eߵ]����\c��qhs)���ͥ@�z��P��trW��fL�yW�(��%3�����}�G˂oٿ˺��܇M$+o��-e]e�6�-�Q�3h��Ș���y�X�%+83{�h��A������������u�{��X�?0��b���<�\l�X�>�+��Upf�9�
�������]�VϹ-��E�>��˱��չ�š��}���Y����BT��[2��L����u�WSd�*���>�T���O���#��[��Wk*�,���s�[��3��p75��eΰ�.B�6 `�)9��;�v��N���yage:���m�q�`a�aĳ���5k���E�d�ff��_lAϊ"������{v�*���d߶4�Y�Y������_���;np�\��9R8��v��N���:<�����#eݕ��m:k:$i:'z%�Z/�N�/�ܕ[�Q�����Ꞧ ϯ��2+��Q��^sV�N�m��̽m�����x���_���}a�	yƳ�<�=��8{�!�?"���1���+�����O�D���H�9�[����5>�g�󾷗��g0�@��;(Z��sG�+X��}wm�B�5���<<�6�����{���$�y�`�lݧ�g�"���1}Z����9�|�/ɼm�I�=���_����������]������w������Ϯ���]�]�o�ͷ?����PK
   -�mVRe��1  ��                  cirkitFile.jsonPK      =   2    